0 0
86 -435
545 -1316
1876 -2808
7343 -7343
-2952 1972
-2759 1143
-2842 565
-2594 0
-2842 -565
-2759 -1143
-2952 -1972
7343 7343
1876 2808
545 1316
86 435
