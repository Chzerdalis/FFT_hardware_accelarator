0 0
0 -33
1 -43
3 -93
5 -112
8 -133
11 -157
16 -190
21 -219
26 -237
34 -277
41 -305
49 -332
58 -366
70 -407
81 -435
94 -473
136 -645
156 -695
131 -553
151 -604
174 -661
291 -1052
198 -685
226 -748
256 -810
284 -862
318 -926
355 -993
402 -1081
474 -1230
1033 -2584
446 -1077
566 -1322
723 -1631
1780 -3887
1753 -3706
1701 -3487
320 -636
548 -1057
693 -1297
805 -1462
926 -1635
1058 -1816
1210 -2019
1385 -2249
1597 -2523
1886 -2899
2316 -3466
3164 -4612
8798 -12492
7615 -10536
6460 -8710
-877 1152
787 -1009
1652 -2064
2473 -3013
3517 -4180
5449 -6317
17214 -19468
12501 -13793
-2198 2366
1931 -2028
4864 -4985
9734 -9734
40208 -39233
10328 -9833
20162 -18730
-14947 13547
4005 -3542
-11908 10272
-7407 6232
-5526 4535
-4171 3338
-2808 2191
-598 455
13020 -9656
-11133 8047
-6584 4637
-5252 3603
-4539 3033
-4062 2643
-3698 2342
-3390 2089
-3118 1869
-2848 1660
-2508 1421
-1964 1081
611 -326
-3722 1931
-663 334
-4068 1985
-1517 717
-4413 2021
-3518 1559
-3199 1371
-3004 1244
-2861 1144
-2731 1053
-2564 953
-1949 697
-3124 1074
-2781 918
-2667 845
-2590 785
-2533 734
-2496 690
-2458 647
-2412 604
-2379 564
-2334 524
-2229 472
-2326 462
-2360 439
-2406 417
-2338 376
-2324 344
-2287 310
-2267 279
-2270 251
-2252 221
-2255 194
-2239 165
-2227 136
-2229 109
-2230 82
-2216 54
-2227 27
-2224 0
-2227 -27
-2216 -54
-2230 -82
-2229 -109
-2227 -136
-2239 -165
-2255 -194
-2252 -221
-2270 -251
-2267 -279
-2287 -310
-2324 -344
-2338 -376
-2406 -417
-2360 -439
-2326 -462
-2229 -472
-2334 -524
-2379 -564
-2412 -604
-2458 -647
-2496 -690
-2533 -734
-2590 -785
-2667 -845
-2781 -918
-3124 -1074
-1949 -697
-2564 -953
-2731 -1053
-2861 -1144
-3004 -1244
-3199 -1371
-3518 -1559
-4413 -2021
-1517 -717
-4068 -1985
-663 -334
-3722 -1931
611 326
-1964 -1081
-2508 -1421
-2848 -1660
-3118 -1869
-3390 -2089
-3698 -2342
-4062 -2643
-4539 -3033
-5252 -3603
-6584 -4637
-11133 -8047
13020 9656
-598 -455
-2808 -2191
-4171 -3338
-5526 -4535
-7407 -6232
-11908 -10272
4005 3542
-14947 -13547
20162 18730
10328 9833
40208 39233
9734 9734
4864 4985
1931 2028
-2198 -2366
12501 13793
17214 19468
5449 6317
3517 4180
2473 3013
1652 2064
787 1009
-877 -1152
6460 8710
7615 10536
8798 12492
3164 4612
2316 3466
1886 2899
1597 2523
1385 2249
1210 2019
1058 1816
926 1635
805 1462
693 1297
548 1057
320 636
1701 3487
1753 3706
1780 3887
723 1631
566 1322
446 1077
1033 2584
474 1230
402 1081
355 993
318 926
284 862
256 810
226 748
198 685
291 1052
174 661
151 604
131 553
156 695
136 645
94 473
81 435
70 407
58 366
49 332
41 305
34 277
26 237
21 219
16 190
11 157
8 133
5 112
3 93
1 43
0 33
