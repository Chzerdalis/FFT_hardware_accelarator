w_real[0] = 9'h0FF; w_imag[0] = 9'h000;
w_real[1] = 9'h0FE; w_imag[1] = 9'h1E7;
w_real[2] = 9'h0FB; w_imag[2] = 9'h1CF;
w_real[3] = 9'h0F4; w_imag[3] = 9'h1B6;
w_real[4] = 9'h0EC; w_imag[4] = 9'h19F;
w_real[5] = 9'h0E1; w_imag[5] = 9'h188;
w_real[6] = 9'h0D4; w_imag[6] = 9'h172;
w_real[7] = 9'h0C5; w_imag[7] = 9'h15E;
w_real[8] = 9'h0B5; w_imag[8] = 9'h14B;
w_real[9] = 9'h0A2; w_imag[9] = 9'h13B;
w_real[10] = 9'h08E; w_imag[10] = 9'h12C;
w_real[11] = 9'h078; w_imag[11] = 9'h11F;
w_real[12] = 9'h061; w_imag[12] = 9'h114;
w_real[13] = 9'h04A; w_imag[13] = 9'h10C;
w_real[14] = 9'h031; w_imag[14] = 9'h105;
w_real[15] = 9'h019; w_imag[15] = 9'h102;
w_real[16] = 9'h000; w_imag[16] = 9'h100;
w_real[17] = 9'h1E7; w_imag[17] = 9'h102;
w_real[18] = 9'h1CF; w_imag[18] = 9'h105;
w_real[19] = 9'h1B6; w_imag[19] = 9'h10C;
w_real[20] = 9'h19F; w_imag[20] = 9'h114;
w_real[21] = 9'h188; w_imag[21] = 9'h11F;
w_real[22] = 9'h172; w_imag[22] = 9'h12C;
w_real[23] = 9'h15E; w_imag[23] = 9'h13B;
w_real[24] = 9'h14B; w_imag[24] = 9'h14B;
w_real[25] = 9'h13B; w_imag[25] = 9'h15E;
w_real[26] = 9'h12C; w_imag[26] = 9'h172;
w_real[27] = 9'h11F; w_imag[27] = 9'h188;
w_real[28] = 9'h114; w_imag[28] = 9'h19F;
w_real[29] = 9'h10C; w_imag[29] = 9'h1B6;
w_real[30] = 9'h105; w_imag[30] = 9'h1CF;
w_real[31] = 9'h102; w_imag[31] = 9'h1E7;
w_real[32] = 9'h100; w_imag[32] = 9'h000;
w_real[33] = 9'h102; w_imag[33] = 9'h019;
w_real[34] = 9'h105; w_imag[34] = 9'h031;
w_real[35] = 9'h10C; w_imag[35] = 9'h04A;
w_real[36] = 9'h114; w_imag[36] = 9'h061;
w_real[37] = 9'h11F; w_imag[37] = 9'h078;
w_real[38] = 9'h12C; w_imag[38] = 9'h08E;
w_real[39] = 9'h13B; w_imag[39] = 9'h0A2;
w_real[40] = 9'h14B; w_imag[40] = 9'h0B5;
w_real[41] = 9'h15E; w_imag[41] = 9'h0C5;
w_real[42] = 9'h172; w_imag[42] = 9'h0D4;
w_real[43] = 9'h188; w_imag[43] = 9'h0E1;
w_real[44] = 9'h19F; w_imag[44] = 9'h0EC;
w_real[45] = 9'h1B6; w_imag[45] = 9'h0F4;
w_real[46] = 9'h1CF; w_imag[46] = 9'h0FB;
w_real[47] = 9'h1E7; w_imag[47] = 9'h0FE;
w_real[48] = 9'h000; w_imag[48] = 9'h0FF;
w_real[49] = 9'h019; w_imag[49] = 9'h0FE;
w_real[50] = 9'h031; w_imag[50] = 9'h0FB;
w_real[51] = 9'h04A; w_imag[51] = 9'h0F4;
w_real[52] = 9'h061; w_imag[52] = 9'h0EC;
w_real[53] = 9'h078; w_imag[53] = 9'h0E1;
w_real[54] = 9'h08E; w_imag[54] = 9'h0D4;
w_real[55] = 9'h0A2; w_imag[55] = 9'h0C5;
w_real[56] = 9'h0B5; w_imag[56] = 9'h0B5;
w_real[57] = 9'h0C5; w_imag[57] = 9'h0A2;
w_real[58] = 9'h0D4; w_imag[58] = 9'h08E;
w_real[59] = 9'h0E1; w_imag[59] = 9'h078;
w_real[60] = 9'h0EC; w_imag[60] = 9'h061;
w_real[61] = 9'h0F4; w_imag[61] = 9'h04A;
w_real[62] = 9'h0FB; w_imag[62] = 9'h031;
w_real[63] = 9'h0FE; w_imag[63] = 9'h019;
