gen_input_real[0] = 18'sd0;
gen_input_real[64] = 18'sd255;
gen_input_real[128] = -18'sd4;
gen_input_real[192] = -18'sd165;
gen_input_real[16] = 18'sd0;
gen_input_real[80] = 18'sd91;
gen_input_real[144] = 18'sd5;
gen_input_real[208] = -18'sd68;
gen_input_real[32] = -18'sd8;
gen_input_real[96] = 18'sd58;
gen_input_real[160] = 18'sd32;
gen_input_real[224] = -18'sd35;
gen_input_real[48] = -18'sd76;
gen_input_real[112] = 18'sd8;
gen_input_real[176] = 18'sd109;
gen_input_real[240] = 18'sd0;
gen_input_real[4] = -18'sd117;
gen_input_real[68] = 18'sd15;
gen_input_real[132] = 18'sd126;
gen_input_real[196] = -18'sd37;
gen_input_real[20] = -18'sd142;
gen_input_real[84] = 18'sd57;
gen_input_real[148] = 18'sd143;
gen_input_real[212] = -18'sd62;
gen_input_real[36] = -18'sd132;
gen_input_real[100] = 18'sd43;
gen_input_real[164] = 18'sd133;
gen_input_real[228] = -18'sd7;
gen_input_real[52] = -18'sd137;
gen_input_real[116] = -18'sd23;
gen_input_real[180] = 18'sd108;
gen_input_real[244] = 18'sd40;
gen_input_real[8] = -18'sd47;
gen_input_real[72] = -18'sd49;
gen_input_real[136] = 18'sd0;
gen_input_real[200] = 18'sd57;
gen_input_real[24] = 18'sd6;
gen_input_real[88] = -18'sd69;
gen_input_real[152] = -18'sd1;
gen_input_real[216] = 18'sd103;
gen_input_real[40] = 18'sd6;
gen_input_real[104] = -18'sd144;
gen_input_real[168] = 18'sd3;
gen_input_real[232] = 18'sd142;
gen_input_real[56] = -18'sd41;
gen_input_real[120] = -18'sd94;
gen_input_real[184] = 18'sd79;
gen_input_real[248] = 18'sd60;
gen_input_real[12] = -18'sd90;
gen_input_real[76] = -18'sd61;
gen_input_real[140] = 18'sd71;
gen_input_real[204] = 18'sd55;
gen_input_real[28] = -18'sd34;
gen_input_real[92] = -18'sd26;
gen_input_real[156] = -18'sd8;
gen_input_real[220] = -18'sd3;
gen_input_real[44] = 18'sd52;
gen_input_real[108] = 18'sd13;
gen_input_real[172] = -18'sd97;
gen_input_real[236] = 18'sd6;
gen_input_real[60] = 18'sd133;
gen_input_real[124] = -18'sd35;
gen_input_real[188] = -18'sd128;
gen_input_real[252] = 18'sd42;
gen_input_real[1] = 18'sd75;
gen_input_real[65] = -18'sd38;
gen_input_real[129] = -18'sd16;
gen_input_real[193] = 18'sd38;
gen_input_real[17] = -18'sd1;
gen_input_real[81] = -18'sd35;
gen_input_real[145] = -18'sd5;
gen_input_real[209] = 18'sd37;
gen_input_real[33] = -18'sd2;
gen_input_real[97] = -18'sd35;
gen_input_real[161] = 18'sd29;
gen_input_real[225] = 18'sd19;
gen_input_real[49] = -18'sd40;
gen_input_real[113] = -18'sd5;
gen_input_real[177] = 18'sd19;
gen_input_real[241] = -18'sd7;
gen_input_real[5] = 18'sd10;
gen_input_real[69] = 18'sd29;
gen_input_real[133] = -18'sd22;
gen_input_real[197] = -18'sd53;
gen_input_real[21] = 18'sd22;
gen_input_real[85] = 18'sd58;
gen_input_real[149] = -18'sd27;
gen_input_real[213] = -18'sd50;
gen_input_real[37] = 18'sd31;
gen_input_real[101] = 18'sd41;
gen_input_real[165] = -18'sd33;
gen_input_real[229] = -18'sd13;
gen_input_real[53] = 18'sd38;
gen_input_real[117] = -18'sd51;
gen_input_real[181] = -18'sd35;
gen_input_real[245] = 18'sd110;
gen_input_real[9] = 18'sd23;
gen_input_real[73] = -18'sd114;
gen_input_real[137] = -18'sd10;
gen_input_real[201] = 18'sd82;
gen_input_real[25] = -18'sd15;
gen_input_real[89] = -18'sd52;
gen_input_real[153] = 18'sd52;
gen_input_real[217] = 18'sd25;
gen_input_real[41] = -18'sd55;
gen_input_real[105] = 18'sd9;
gen_input_real[169] = 18'sd4;
gen_input_real[233] = -18'sd52;
gen_input_real[57] = 18'sd48;
gen_input_real[121] = 18'sd79;
gen_input_real[185] = -18'sd50;
gen_input_real[249] = -18'sd73;
gen_input_real[13] = 18'sd23;
gen_input_real[77] = 18'sd45;
gen_input_real[141] = -18'sd32;
gen_input_real[205] = -18'sd6;
gen_input_real[29] = 18'sd80;
gen_input_real[93] = -18'sd39;
gen_input_real[157] = -18'sd105;
gen_input_real[221] = 18'sd62;
gen_input_real[45] = 18'sd80;
gen_input_real[109] = -18'sd43;
gen_input_real[173] = -18'sd44;
gen_input_real[237] = 18'sd13;
gen_input_real[61] = 18'sd31;
gen_input_real[125] = 18'sd0;
gen_input_real[189] = -18'sd28;
gen_input_real[253] = -18'sd13;
gen_input_real[2] = 18'sd13;
gen_input_real[66] = 18'sd28;
gen_input_real[130] = 18'sd0;
gen_input_real[194] = -18'sd31;
gen_input_real[18] = -18'sd13;
gen_input_real[82] = 18'sd44;
gen_input_real[146] = 18'sd43;
gen_input_real[210] = -18'sd80;
gen_input_real[34] = -18'sd62;
gen_input_real[98] = 18'sd105;
gen_input_real[162] = 18'sd39;
gen_input_real[226] = -18'sd80;
gen_input_real[50] = 18'sd6;
gen_input_real[114] = 18'sd32;
gen_input_real[178] = -18'sd45;
gen_input_real[242] = -18'sd23;
gen_input_real[6] = 18'sd73;
gen_input_real[70] = 18'sd50;
gen_input_real[134] = -18'sd79;
gen_input_real[198] = -18'sd48;
gen_input_real[22] = 18'sd52;
gen_input_real[86] = -18'sd4;
gen_input_real[150] = -18'sd9;
gen_input_real[214] = 18'sd55;
gen_input_real[38] = -18'sd25;
gen_input_real[102] = -18'sd52;
gen_input_real[166] = 18'sd52;
gen_input_real[230] = 18'sd15;
gen_input_real[54] = -18'sd82;
gen_input_real[118] = 18'sd10;
gen_input_real[182] = 18'sd114;
gen_input_real[246] = -18'sd23;
gen_input_real[10] = -18'sd110;
gen_input_real[74] = 18'sd35;
gen_input_real[138] = 18'sd51;
gen_input_real[202] = -18'sd38;
gen_input_real[26] = 18'sd13;
gen_input_real[90] = 18'sd33;
gen_input_real[154] = -18'sd41;
gen_input_real[218] = -18'sd31;
gen_input_real[42] = 18'sd50;
gen_input_real[106] = 18'sd27;
gen_input_real[170] = -18'sd58;
gen_input_real[234] = -18'sd22;
gen_input_real[58] = 18'sd53;
gen_input_real[122] = 18'sd22;
gen_input_real[186] = -18'sd29;
gen_input_real[250] = -18'sd10;
gen_input_real[14] = 18'sd7;
gen_input_real[78] = -18'sd19;
gen_input_real[142] = 18'sd5;
gen_input_real[206] = 18'sd40;
gen_input_real[30] = -18'sd19;
gen_input_real[94] = -18'sd29;
gen_input_real[158] = 18'sd35;
gen_input_real[222] = 18'sd2;
gen_input_real[46] = -18'sd37;
gen_input_real[110] = 18'sd5;
gen_input_real[174] = 18'sd35;
gen_input_real[238] = 18'sd1;
gen_input_real[62] = -18'sd38;
gen_input_real[126] = 18'sd16;
gen_input_real[190] = 18'sd38;
gen_input_real[254] = -18'sd75;
gen_input_real[3] = -18'sd42;
gen_input_real[67] = 18'sd128;
gen_input_real[131] = 18'sd35;
gen_input_real[195] = -18'sd133;
gen_input_real[19] = -18'sd6;
gen_input_real[83] = 18'sd97;
gen_input_real[147] = -18'sd13;
gen_input_real[211] = -18'sd52;
gen_input_real[35] = 18'sd3;
gen_input_real[99] = 18'sd8;
gen_input_real[163] = 18'sd26;
gen_input_real[227] = 18'sd34;
gen_input_real[51] = -18'sd55;
gen_input_real[115] = -18'sd71;
gen_input_real[179] = 18'sd61;
gen_input_real[243] = 18'sd90;
gen_input_real[7] = -18'sd60;
gen_input_real[71] = -18'sd79;
gen_input_real[135] = 18'sd94;
gen_input_real[199] = 18'sd41;
gen_input_real[23] = -18'sd142;
gen_input_real[87] = -18'sd3;
gen_input_real[151] = 18'sd144;
gen_input_real[215] = -18'sd6;
gen_input_real[39] = -18'sd103;
gen_input_real[103] = 18'sd1;
gen_input_real[167] = 18'sd69;
gen_input_real[231] = -18'sd6;
gen_input_real[55] = -18'sd57;
gen_input_real[119] = 18'sd0;
gen_input_real[183] = 18'sd49;
gen_input_real[247] = 18'sd47;
gen_input_real[11] = -18'sd40;
gen_input_real[75] = -18'sd108;
gen_input_real[139] = 18'sd23;
gen_input_real[203] = 18'sd137;
gen_input_real[27] = 18'sd7;
gen_input_real[91] = -18'sd133;
gen_input_real[155] = -18'sd43;
gen_input_real[219] = 18'sd132;
gen_input_real[43] = 18'sd62;
gen_input_real[107] = -18'sd143;
gen_input_real[171] = -18'sd57;
gen_input_real[235] = 18'sd142;
gen_input_real[59] = 18'sd37;
gen_input_real[123] = -18'sd126;
gen_input_real[187] = -18'sd15;
gen_input_real[251] = 18'sd117;
gen_input_real[15] = 18'sd0;
gen_input_real[79] = -18'sd109;
gen_input_real[143] = -18'sd8;
gen_input_real[207] = 18'sd76;
gen_input_real[31] = 18'sd35;
gen_input_real[95] = -18'sd32;
gen_input_real[159] = -18'sd58;
gen_input_real[223] = 18'sd8;
gen_input_real[47] = 18'sd68;
gen_input_real[111] = -18'sd5;
gen_input_real[175] = -18'sd91;
gen_input_real[239] = 18'sd0;
gen_input_real[63] = 18'sd165;
gen_input_real[127] = 18'sd4;
gen_input_real[191] = -18'sd255;
gen_input_real[255] = 18'sd0;
