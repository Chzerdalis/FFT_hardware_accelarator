0 0
5 -432
21 -868
47 -1301
85 -1730
134 -2188
193 -2617
264 -3069
344 -3499
440 -3970
547 -4436
667 -4916
800 -5399
950 -5906
1116 -6432
1300 -6984
1515 -7618
2186 -10329
2499 -11129
2103 -8856
2423 -9675
2787 -10577
4659 -16837
3166 -10917
3631 -11971
4078 -12873
4556 -13793
5090 -14796
5706 -15948
6468 -17402
7609 -19726
16532 -41341
7121 -17193
9100 -21229
11551 -26059
28465 -62146
28068 -59345
27248 -55828
5042 -10017
8838 -17034
11039 -20653
12946 -23522
14858 -26229
16932 -29051
19279 -32165
22070 -35818
25536 -40326
30178 -46387
37153 -55603
50679 -73867
140874 -200026
121963 -168738
103431 -139460
-14053 18470
12500 -16017
26458 -33058
39510 -48144
56304 -66915
87095 -100968
275782 -311886
200339 -221041
-35281 37979
30878 -32432
77720 -79651
155961 -155961
644199 -628579
165440 -157512
322955 -300009
-239484 217056
64157 -56730
-190789 164576
-118777 99942
-88324 72485
-66722 53401
-45071 35174
-9596 7301
208622 -154724
-178346 128908
-105483 74289
-84032 57652
-72648 48542
-65024 42303
-59236 37510
-54403 33522
-50006 29972
-45547 26545
-40204 22775
-31440 17304
9862 -5271
-59793 31023
-10724 5398
-65117 31782
-24384 11532
-70699 32382
-56213 24917
-51204 21949
-48155 19946
-45809 18319
-43675 16847
-40988 15236
-31257 11184
-50156 17254
-44516 14706
-42667 13517
-41516 12593
-40633 11783
-39910 11044
-39276 10352
-38670 9686
-38087 9045
-37394 8397
-35712 7560
-37219 7403
-37694 7018
-38352 6654
-37399 6017
-36970 5484
-36644 4976
-36292 4476
-36424 4039
-36164 3561
-36000 3100
-35872 2646
-35764 2197
-35678 1752
-35641 1312
-35595 873
-35568 436
-35550 0
-35568 -436
-35595 -873
-35641 -1312
-35678 -1752
-35764 -2197
-35872 -2646
-36000 -3100
-36164 -3561
-36424 -4039
-36292 -4476
-36644 -4976
-36970 -5484
-37399 -6017
-38352 -6654
-37694 -7018
-37219 -7403
-35712 -7560
-37394 -8397
-38087 -9045
-38670 -9686
-39276 -10352
-39910 -11044
-40633 -11783
-41516 -12593
-42667 -13517
-44516 -14706
-50156 -17254
-31257 -11184
-40988 -15236
-43675 -16847
-45809 -18319
-48155 -19946
-51204 -21949
-56213 -24917
-70699 -32382
-24384 -11532
-65117 -31782
-10724 -5398
-59793 -31023
9862 5271
-31440 -17304
-40204 -22775
-45547 -26545
-50006 -29972
-54403 -33522
-59236 -37510
-65024 -42303
-72648 -48542
-84032 -57652
-105483 -74289
-178346 -128908
208622 154724
-9596 -7301
-45071 -35174
-66722 -53401
-88324 -72485
-118777 -99942
-190789 -164576
64157 56730
-239484 -217056
322955 300009
165440 157512
644199 628579
155961 155961
77720 79651
30878 32432
-35281 -37979
200339 221041
275782 311886
87095 100968
56304 66915
39510 48144
26458 33058
12500 16017
-14053 -18470
103431 139460
121963 168738
140874 200026
50679 73867
37153 55603
30178 46387
25536 40326
22070 35818
19279 32165
16932 29051
14858 26229
12946 23522
11039 20653
8838 17034
5042 10017
27248 55828
28068 59345
28465 62146
11551 26059
9100 21229
7121 17193
16532 41341
7609 19726
6468 17402
5706 15948
5090 14796
4556 13793
4078 12873
3631 11971
3166 10917
4659 16837
2787 10577
2423 9675
2103 8856
2499 11129
2186 10329
1515 7618
1300 6984
1116 6432
950 5906
800 5399
667 4916
547 4436
440 3970
344 3499
264 3069
193 2617
134 2188
85 1730
47 1301
21 868
5 432
