gen_input_real[0] = 16'sd0;
gen_input_real[64] = 16'sd127;
gen_input_real[128] = -16'sd2;
gen_input_real[192] = -16'sd100;
gen_input_real[16] = 16'sd6;
gen_input_real[80] = 16'sd75;
gen_input_real[144] = -16'sd10;
gen_input_real[208] = -16'sd61;
gen_input_real[32] = 16'sd15;
gen_input_real[96] = 16'sd50;
gen_input_real[160] = -16'sd21;
gen_input_real[224] = -16'sd35;
gen_input_real[48] = 16'sd30;
gen_input_real[112] = 16'sd23;
gen_input_real[176] = -16'sd36;
gen_input_real[240] = -16'sd27;
gen_input_real[4] = 16'sd36;
gen_input_real[68] = 16'sd40;
gen_input_real[132] = -16'sd31;
gen_input_real[196] = -16'sd43;
gen_input_real[20] = 16'sd30;
gen_input_real[84] = 16'sd30;
gen_input_real[148] = -16'sd35;
gen_input_real[212] = -16'sd6;
gen_input_real[36] = 16'sd38;
gen_input_real[100] = -16'sd15;
gen_input_real[164] = -16'sd38;
gen_input_real[228] = 16'sd31;
gen_input_real[52] = 16'sd39;
gen_input_real[116] = -16'sd45;
gen_input_real[180] = -16'sd42;
gen_input_real[244] = 16'sd55;
gen_input_real[8] = 16'sd46;
gen_input_real[72] = -16'sd54;
gen_input_real[136] = -16'sd47;
gen_input_real[200] = 16'sd38;
gen_input_real[24] = 16'sd42;
gen_input_real[88] = -16'sd18;
gen_input_real[152] = -16'sd35;
gen_input_real[216] = 16'sd7;
gen_input_real[40] = 16'sd30;
gen_input_real[104] = -16'sd3;
gen_input_real[168] = -16'sd34;
gen_input_real[232] = 16'sd3;
gen_input_real[56] = 16'sd38;
gen_input_real[120] = -16'sd8;
gen_input_real[184] = -16'sd37;
gen_input_real[248] = 16'sd16;
gen_input_real[12] = 16'sd33;
gen_input_real[76] = -16'sd26;
gen_input_real[140] = -16'sd33;
gen_input_real[204] = 16'sd28;
gen_input_real[28] = 16'sd32;
gen_input_real[92] = -16'sd19;
gen_input_real[156] = -16'sd26;
gen_input_real[220] = 16'sd6;
gen_input_real[44] = 16'sd14;
gen_input_real[108] = 16'sd1;
gen_input_real[172] = -16'sd6;
gen_input_real[236] = -16'sd7;
gen_input_real[60] = 16'sd2;
gen_input_real[124] = 16'sd15;
gen_input_real[188] = -16'sd1;
gen_input_real[252] = -16'sd17;
gen_input_real[1] = 16'sd3;
gen_input_real[65] = 16'sd7;
gen_input_real[129] = -16'sd4;
gen_input_real[193] = 16'sd7;
gen_input_real[17] = 16'sd2;
gen_input_real[81] = -16'sd17;
gen_input_real[145] = 16'sd1;
gen_input_real[209] = 16'sd21;
gen_input_real[33] = -16'sd6;
gen_input_real[97] = -16'sd23;
gen_input_real[161] = 16'sd13;
gen_input_real[225] = 16'sd21;
gen_input_real[49] = -16'sd19;
gen_input_real[113] = -16'sd14;
gen_input_real[177] = 16'sd22;
gen_input_real[241] = 16'sd8;
gen_input_real[5] = -16'sd20;
gen_input_real[69] = -16'sd3;
gen_input_real[133] = 16'sd13;
gen_input_real[197] = -16'sd1;
gen_input_real[21] = -16'sd2;
gen_input_real[85] = 16'sd1;
gen_input_real[149] = -16'sd7;
gen_input_real[213] = 16'sd4;
gen_input_real[37] = 16'sd14;
gen_input_real[101] = -16'sd12;
gen_input_real[165] = -16'sd17;
gen_input_real[229] = 16'sd18;
gen_input_real[53] = 16'sd16;
gen_input_real[117] = -16'sd21;
gen_input_real[181] = -16'sd11;
gen_input_real[245] = 16'sd21;
gen_input_real[9] = 16'sd8;
gen_input_real[73] = -16'sd18;
gen_input_real[137] = -16'sd11;
gen_input_real[201] = 16'sd16;
gen_input_real[25] = 16'sd17;
gen_input_real[89] = -16'sd15;
gen_input_real[153] = -16'sd21;
gen_input_real[217] = 16'sd11;
gen_input_real[41] = 16'sd26;
gen_input_real[105] = -16'sd7;
gen_input_real[169] = -16'sd34;
gen_input_real[233] = 16'sd11;
gen_input_real[57] = 16'sd38;
gen_input_real[121] = -16'sd24;
gen_input_real[185] = -16'sd32;
gen_input_real[249] = 16'sd39;
gen_input_real[13] = 16'sd18;
gen_input_real[77] = -16'sd46;
gen_input_real[141] = -16'sd2;
gen_input_real[205] = 16'sd46;
gen_input_real[29] = -16'sd9;
gen_input_real[93] = -16'sd47;
gen_input_real[157] = 16'sd16;
gen_input_real[221] = 16'sd50;
gen_input_real[45] = -16'sd18;
gen_input_real[109] = -16'sd47;
gen_input_real[173] = 16'sd22;
gen_input_real[237] = 16'sd34;
gen_input_real[61] = -16'sd26;
gen_input_real[125] = -16'sd19;
gen_input_real[189] = 16'sd22;
gen_input_real[253] = 16'sd16;
gen_input_real[2] = -16'sd16;
gen_input_real[66] = -16'sd22;
gen_input_real[130] = 16'sd19;
gen_input_real[194] = 16'sd26;
gen_input_real[18] = -16'sd34;
gen_input_real[82] = -16'sd22;
gen_input_real[146] = 16'sd47;
gen_input_real[210] = 16'sd18;
gen_input_real[34] = -16'sd50;
gen_input_real[98] = -16'sd16;
gen_input_real[162] = 16'sd47;
gen_input_real[226] = 16'sd9;
gen_input_real[50] = -16'sd46;
gen_input_real[114] = 16'sd2;
gen_input_real[178] = 16'sd46;
gen_input_real[242] = -16'sd18;
gen_input_real[6] = -16'sd39;
gen_input_real[70] = 16'sd32;
gen_input_real[134] = 16'sd24;
gen_input_real[198] = -16'sd38;
gen_input_real[22] = -16'sd11;
gen_input_real[86] = 16'sd34;
gen_input_real[150] = 16'sd7;
gen_input_real[214] = -16'sd26;
gen_input_real[38] = -16'sd11;
gen_input_real[102] = 16'sd21;
gen_input_real[166] = 16'sd15;
gen_input_real[230] = -16'sd17;
gen_input_real[54] = -16'sd16;
gen_input_real[118] = 16'sd11;
gen_input_real[182] = 16'sd18;
gen_input_real[246] = -16'sd8;
gen_input_real[10] = -16'sd21;
gen_input_real[74] = 16'sd11;
gen_input_real[138] = 16'sd21;
gen_input_real[202] = -16'sd16;
gen_input_real[26] = -16'sd18;
gen_input_real[90] = 16'sd17;
gen_input_real[154] = 16'sd12;
gen_input_real[218] = -16'sd14;
gen_input_real[42] = -16'sd4;
gen_input_real[106] = 16'sd7;
gen_input_real[170] = -16'sd1;
gen_input_real[234] = 16'sd2;
gen_input_real[58] = 16'sd1;
gen_input_real[122] = -16'sd13;
gen_input_real[186] = 16'sd3;
gen_input_real[250] = 16'sd20;
gen_input_real[14] = -16'sd8;
gen_input_real[78] = -16'sd22;
gen_input_real[142] = 16'sd14;
gen_input_real[206] = 16'sd19;
gen_input_real[30] = -16'sd21;
gen_input_real[94] = -16'sd13;
gen_input_real[158] = 16'sd23;
gen_input_real[222] = 16'sd6;
gen_input_real[46] = -16'sd21;
gen_input_real[110] = -16'sd1;
gen_input_real[174] = 16'sd17;
gen_input_real[238] = -16'sd2;
gen_input_real[62] = -16'sd7;
gen_input_real[126] = 16'sd4;
gen_input_real[190] = -16'sd7;
gen_input_real[254] = -16'sd3;
gen_input_real[3] = 16'sd17;
gen_input_real[67] = 16'sd1;
gen_input_real[131] = -16'sd15;
gen_input_real[195] = -16'sd2;
gen_input_real[19] = 16'sd7;
gen_input_real[83] = 16'sd6;
gen_input_real[147] = -16'sd1;
gen_input_real[211] = -16'sd14;
gen_input_real[35] = -16'sd6;
gen_input_real[99] = 16'sd26;
gen_input_real[163] = 16'sd19;
gen_input_real[227] = -16'sd32;
gen_input_real[51] = -16'sd28;
gen_input_real[115] = 16'sd33;
gen_input_real[179] = 16'sd26;
gen_input_real[243] = -16'sd33;
gen_input_real[7] = -16'sd16;
gen_input_real[71] = 16'sd37;
gen_input_real[135] = 16'sd8;
gen_input_real[199] = -16'sd38;
gen_input_real[23] = -16'sd3;
gen_input_real[87] = 16'sd34;
gen_input_real[151] = 16'sd3;
gen_input_real[215] = -16'sd30;
gen_input_real[39] = -16'sd7;
gen_input_real[103] = 16'sd35;
gen_input_real[167] = 16'sd18;
gen_input_real[231] = -16'sd42;
gen_input_real[55] = -16'sd38;
gen_input_real[119] = 16'sd47;
gen_input_real[183] = 16'sd54;
gen_input_real[247] = -16'sd46;
gen_input_real[11] = -16'sd55;
gen_input_real[75] = 16'sd42;
gen_input_real[139] = 16'sd45;
gen_input_real[203] = -16'sd39;
gen_input_real[27] = -16'sd31;
gen_input_real[91] = 16'sd38;
gen_input_real[155] = 16'sd15;
gen_input_real[219] = -16'sd38;
gen_input_real[43] = 16'sd6;
gen_input_real[107] = 16'sd35;
gen_input_real[171] = -16'sd30;
gen_input_real[235] = -16'sd30;
gen_input_real[59] = 16'sd43;
gen_input_real[123] = 16'sd31;
gen_input_real[187] = -16'sd40;
gen_input_real[251] = -16'sd36;
gen_input_real[15] = 16'sd27;
gen_input_real[79] = 16'sd36;
gen_input_real[143] = -16'sd23;
gen_input_real[207] = -16'sd30;
gen_input_real[31] = 16'sd35;
gen_input_real[95] = 16'sd21;
gen_input_real[159] = -16'sd50;
gen_input_real[223] = -16'sd15;
gen_input_real[47] = 16'sd61;
gen_input_real[111] = 16'sd10;
gen_input_real[175] = -16'sd75;
gen_input_real[239] = -16'sd6;
gen_input_real[63] = 16'sd100;
gen_input_real[127] = 16'sd2;
gen_input_real[191] = -16'sd127;
gen_input_real[255] = 16'sd0;
