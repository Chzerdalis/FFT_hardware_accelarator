0 0
0 5
0 6
0 0
0 8
0 2
0 5
0 -14
0 4
0 16
0 5
0 -6
0 14
0 -15
0 -14
0 0
0 -2
0 -1
0 -4
0 -9
0 -4
0 14
0 -8
-1 14
0 -3
0 -12
1 -14
1 -14
2 -23
0 -2
0 1
0 3
0 -5
0 0
4 -38
2 -24
1 -15
1 -14
0 1
3 -27
3 -27
3 -25
4 -34
2 -15
3 -23
1 -12
1 -10
4 -31
2 -17
3 -25
2 -18
2 -14
5 -36
2 -17
4 -25
5 -32
6 -36
5 -29
1 -10
7 -39
3 -16
14 -76
9 -50
2 -14
4 -24
7 -39
7 -35
8 -40
8 -38
7 -36
8 -39
6 -28
13 -60
21 -94
7 -34
6 -29
4 -19
7 -32
9 -40
9 -38
11 -44
18 -72
9 -37
8 -33
9 -37
11 -44
13 -50
18 -69
9 -35
18 -66
8 -29
15 -55
18 -64
12 -44
12 -41
10 -35
19 -63
16 -52
20 -65
22 -71
22 -71
22 -68
15 -48
26 -80
24 -75
24 -73
29 -86
32 -95
142 -413
18 -53
25 -72
156 -442
-1 3
11 -32
15 -42
28 -77
24 -66
26 -70
33 -87
221 -579
2 -7
16 -41
16 -40
19 -49
24 -62
30 -76
24 -60
27 -68
21 -52
30 -73
38 -90
33 -79
39 -92
26 -60
36 -84
39 -89
44 -100
44 -98
41 -92
54 -120
54 -119
63 -136
73 -157
97 -207
529 -1120
-35 74
5 -10
19 -40
30 -62
29 -60
45 -92
43 -86
40 -79
59 -116
62 -121
51 -99
53 -102
69 -132
73 -139
79 -148
91 -171
101 -187
121 -223
191 -349
980 -1780
-127 230
-25 45
21 -38
30 -54
38 -67
46 -80
62 -107
53 -91
65 -111
71 -120
54 -91
82 -137
83 -138
86 -142
90 -148
96 -156
104 -167
121 -194
122 -195
148 -234
186 -292
225 -351
354 -548
1844 -2834
-305 467
-86 130
-1 2
39 -58
65 -96
85 -126
96 -141
109 -160
149 -216
200 -288
276 -395
446 -634
2486 -3507
-522 732
-193 269
-74 102
-41 57
-14 19
4 -6
48 -65
47 -63
56 -75
74 -98
90 -119
95 -125
116 -151
116 -150
131 -168
166 -211
200 -253
217 -273
240 -300
273 -339
370 -456
493 -605
821 -1000
4213 -5102
-1059 1275
-387 463
-196 233
-113 134
-72 84
-9 10
-1 1
30 -34
62 -71
91 -104
105 -119
137 -154
165 -184
190 -211
204 -226
214 -235
238 -260
288 -312
350 -377
383 -410
455 -484
519 -548
629 -660
794 -829
1095 -1136
1798 -1854
7500 -7686
-1461 1489
488 -494
6735 -6777
-2869 2869
-1368 1359
-914 903
-703 690
-562 549
-443 429
-376 363
-321 308
-269 256
-235 222
-205 193
-151 142
-123 114
-67 62
-4 3
52 -47
120 -109
263 -237
475 -425
1009 -898
5440 -4810
-2239 1968
-1035 904
-685 595
-580 500
-475 407
-412 351
-343 290
-339 285
-293 245
-268 222
-240 198
-221 182
-203 165
-186 151
-154 124
-171 137
-157 124
-132 104
-137 107
-96 75
-98 76
-66 50
-73 56
-34 26
-39 29
3 -2
42 -31
115 -85
174 -128
327 -239
649 -472
3154 -2279
-1551 1113
-700 500
-455 323
-379 267
-303 212
-270 187
-227 156
-208 142
-198 135
-160 108
-134 90
-129 86
-108 71
-110 72
-106 69
-96 62
-47 30
-56 36
-2 1
-12 8
32 -20
54 -33
115 -71
201 -124
421 -257
1924 -1169
-966 583
-376 225
-200 119
-83 49
-26 15
108 -63
300 -174
1598 -918
-789 450
-246 139
74 -41
1257 -702
-900 499
-394 217
-166 90
66 -35
1148 -618
-688 368
695 -368
-1106 582
-657 343
-511 265
-452 233
-373 190
-353 179
-329 165
-313 156
-298 147
-259 127
-235 115
-236 114
-213 102
-191 91
-189 89
-115 53
-40 18
564 -260
-672 308
-418 190
-338 152
-283 126
-278 123
-259 114
-246 107
-222 96
-218 93
-215 91
-208 88
-194 81
-197 81
-208 85
-179 72
-157 63
-141 56
-134 53
-72 28
262 -102
-436 168
-267 102
-194 73
-123 46
112 -41
-446 164
-321 117
-238 86
-220 79
-228 80
-215 75
-207 72
-191 65
-187 63
-173 58
-144 48
40 -13
-358 117
-271 87
-241 77
-225 71
-192 60
-207 64
-192 59
-192 58
-186 55
-193 57
-154 45
-70 20
-280 80
-222 63
-225 63
-191 52
-228 62
-183 49
-178 47
-169 44
-189 49
-176 45
-192 48
-165 41
-166 41
-172 42
-190 45
-169 40
-176 41
-190 44
-159 36
-163 36
-165 36
-181 39
-191 41
-160 33
-162 33
-167 34
-160 32
-182 36
-163 31
-174 33
-168 31
-145 27
-169 31
-157 28
-167 29
-154 26
-159 27
-158 26
-159 26
-162 26
-177 27
-151 23
-165 25
-173 25
-156 22
-163 23
-146 20
-150 20
-144 19
-148 19
-175 22
-160 19
-172 20
-159 18
-167 19
-145 16
-159 17
-145 15
-165 16
-165 16
-163 15
-149 13
-176 15
-154 13
-172 14
-158 12
-150 11
-161 11
-158 11
-144 9
-170 11
-140 8
-165 9
-127 7
-153 8
-165 8
-146 6
-161 6
-168 6
-152 5
-162 5
-150 4
-144 3
-156 3
-161 3
-142 2
-176 2
-164 2
-163 1
-177 1
-181 0
-158 0
-181 0
-177 -1
-163 -1
-164 -2
-176 -2
-142 -2
-161 -3
-156 -3
-144 -3
-150 -4
-162 -5
-152 -5
-168 -6
-161 -6
-146 -6
-165 -8
-153 -8
-127 -7
-165 -9
-140 -8
-170 -11
-144 -9
-158 -11
-161 -11
-150 -11
-158 -12
-172 -14
-154 -13
-176 -15
-149 -13
-163 -15
-165 -16
-165 -16
-145 -15
-159 -17
-145 -16
-167 -19
-159 -18
-172 -20
-160 -19
-175 -22
-148 -19
-144 -19
-150 -20
-146 -20
-163 -23
-156 -22
-173 -25
-165 -25
-151 -23
-177 -27
-162 -26
-159 -26
-158 -26
-159 -27
-154 -26
-167 -29
-157 -28
-169 -31
-145 -27
-168 -31
-174 -33
-163 -31
-182 -36
-160 -32
-167 -34
-162 -33
-160 -33
-191 -41
-181 -39
-165 -36
-163 -36
-159 -36
-190 -44
-176 -41
-169 -40
-190 -45
-172 -42
-166 -41
-165 -41
-192 -48
-176 -45
-189 -49
-169 -44
-178 -47
-183 -49
-228 -62
-191 -52
-225 -63
-222 -63
-280 -80
-70 -20
-154 -45
-193 -57
-186 -55
-192 -58
-192 -59
-207 -64
-192 -60
-225 -71
-241 -77
-271 -87
-358 -117
40 13
-144 -48
-173 -58
-187 -63
-191 -65
-207 -72
-215 -75
-228 -80
-220 -79
-238 -86
-321 -117
-446 -164
112 41
-123 -46
-194 -73
-267 -102
-436 -168
262 102
-72 -28
-134 -53
-141 -56
-157 -63
-179 -72
-208 -85
-197 -81
-194 -81
-208 -88
-215 -91
-218 -93
-222 -96
-246 -107
-259 -114
-278 -123
-283 -126
-338 -152
-418 -190
-672 -308
564 260
-40 -18
-115 -53
-189 -89
-191 -91
-213 -102
-236 -114
-235 -115
-259 -127
-298 -147
-313 -156
-329 -165
-353 -179
-373 -190
-452 -233
-511 -265
-657 -343
-1106 -582
695 368
-688 -368
1148 618
66 35
-166 -90
-394 -217
-900 -499
1257 702
74 41
-246 -139
-789 -450
1598 918
300 174
108 63
-26 -15
-83 -49
-200 -119
-376 -225
-966 -583
1924 1169
421 257
201 124
115 71
54 33
32 20
-12 -8
-2 -1
-56 -36
-47 -30
-96 -62
-106 -69
-110 -72
-108 -71
-129 -86
-134 -90
-160 -108
-198 -135
-208 -142
-227 -156
-270 -187
-303 -212
-379 -267
-455 -323
-700 -500
-1551 -1113
3154 2279
649 472
327 239
174 128
115 85
42 31
3 2
-39 -29
-34 -26
-73 -56
-66 -50
-98 -76
-96 -75
-137 -107
-132 -104
-157 -124
-171 -137
-154 -124
-186 -151
-203 -165
-221 -182
-240 -198
-268 -222
-293 -245
-339 -285
-343 -290
-412 -351
-475 -407
-580 -500
-685 -595
-1035 -904
-2239 -1968
5440 4810
1009 898
475 425
263 237
120 109
52 47
-4 -3
-67 -62
-123 -114
-151 -142
-205 -193
-235 -222
-269 -256
-321 -308
-376 -363
-443 -429
-562 -549
-703 -690
-914 -903
-1368 -1359
-2869 -2869
6735 6777
488 494
-1461 -1489
7500 7686
1798 1854
1095 1136
794 829
629 660
519 548
455 484
383 410
350 377
288 312
238 260
214 235
204 226
190 211
165 184
137 154
105 119
91 104
62 71
30 34
-1 -1
-9 -10
-72 -84
-113 -134
-196 -233
-387 -463
-1059 -1275
4213 5102
821 1000
493 605
370 456
273 339
240 300
217 273
200 253
166 211
131 168
116 150
116 151
95 125
90 119
74 98
56 75
47 63
48 65
4 6
-14 -19
-41 -57
-74 -102
-193 -269
-522 -732
2486 3507
446 634
276 395
200 288
149 216
109 160
96 141
85 126
65 96
39 58
-1 -2
-86 -130
-305 -467
1844 2834
354 548
225 351
186 292
148 234
122 195
121 194
104 167
96 156
90 148
86 142
83 138
82 137
54 91
71 120
65 111
53 91
62 107
46 80
38 67
30 54
21 38
-25 -45
-127 -230
980 1780
191 349
121 223
101 187
91 171
79 148
73 139
69 132
53 102
51 99
62 121
59 116
40 79
43 86
45 92
29 60
30 62
19 40
5 10
-35 -74
529 1120
97 207
73 157
63 136
54 119
54 120
41 92
44 98
44 100
39 89
36 84
26 60
39 92
33 79
38 90
30 73
21 52
27 68
24 60
30 76
24 62
19 49
16 40
16 41
2 7
221 579
33 87
26 70
24 66
28 77
15 42
11 32
-1 -3
156 442
25 72
18 53
142 413
32 95
29 86
24 73
24 75
26 80
15 48
22 68
22 71
22 71
20 65
16 52
19 63
10 35
12 41
12 44
18 64
15 55
8 29
18 66
9 35
18 69
13 50
11 44
9 37
8 33
9 37
18 72
11 44
9 38
9 40
7 32
4 19
6 29
7 34
21 94
13 60
6 28
8 39
7 36
8 38
8 40
7 35
7 39
4 24
2 14
9 50
14 76
3 16
7 39
1 10
5 29
6 36
5 32
4 25
2 17
5 36
2 14
2 18
3 25
2 17
4 31
1 10
1 12
3 23
2 15
4 34
3 25
3 27
3 27
0 -1
1 14
1 15
2 24
4 38
0 0
0 5
0 -3
0 -1
0 2
2 23
1 14
1 14
0 12
0 3
-1 -14
0 8
0 -14
0 4
0 9
0 4
0 1
0 2
0 0
0 14
0 15
0 -14
0 6
0 -5
0 -16
0 -4
0 14
0 -5
0 -2
0 -8
0 0
0 -6
0 -5
