0 0
5 -115
23 -234
52 -356
118 -597
160 -638
347 -1144
339 -949
510 -1232
769 -1627
1233 -2308
3709 -6189
5679 -8500
834 -1124
7937 -9671
4222 -4658
5385 -5385
6444 -5841
-2565 2105
-5294 3926
-3443 2300
-2571 1541
-1194 638
-1464 692
-2548 1055
-3269 1169
-2673 811
-2411 604
-2391 475
-2310 342
-2274 224
-2242 110
-2238 0
-2242 -110
-2274 -224
-2310 -342
-2391 -475
-2411 -604
-2673 -811
-3269 -1169
-2548 -1055
-1464 -692
-1194 -638
-2571 -1541
-3443 -2300
-5294 -3926
-2565 -2105
6444 5841
5385 5385
4222 4658
7937 9671
834 1124
5679 8500
3709 6189
1233 2308
769 1627
510 1232
339 949
347 1144
160 638
118 597
52 356
23 234
5 115
