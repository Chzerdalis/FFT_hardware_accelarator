w_real[0] = 8'h7F; w_imag[0] = 8'h00;
w_real[1] = 8'h7F; w_imag[1] = 8'h00;
w_real[2] = 8'h7F; w_imag[2] = 8'hFF;
w_real[3] = 8'h7F; w_imag[3] = 8'hFE;
w_real[4] = 8'h7F; w_imag[4] = 8'hFD;
w_real[5] = 8'h7F; w_imag[5] = 8'hFD;
w_real[6] = 8'h7F; w_imag[6] = 8'hFC;
w_real[7] = 8'h7F; w_imag[7] = 8'hFB;
w_real[8] = 8'h7F; w_imag[8] = 8'hFA;
w_real[9] = 8'h7F; w_imag[9] = 8'hF9;
w_real[10] = 8'h7F; w_imag[10] = 8'hF9;
w_real[11] = 8'h7F; w_imag[11] = 8'hF8;
w_real[12] = 8'h7F; w_imag[12] = 8'hF7;
w_real[13] = 8'h7F; w_imag[13] = 8'hF6;
w_real[14] = 8'h7F; w_imag[14] = 8'hF6;
w_real[15] = 8'h7F; w_imag[15] = 8'hF5;
w_real[16] = 8'h7F; w_imag[16] = 8'hF4;
w_real[17] = 8'h7F; w_imag[17] = 8'hF3;
w_real[18] = 8'h7F; w_imag[18] = 8'hF2;
w_real[19] = 8'h7F; w_imag[19] = 8'hF2;
w_real[20] = 8'h7F; w_imag[20] = 8'hF1;
w_real[21] = 8'h7E; w_imag[21] = 8'hF0;
w_real[22] = 8'h7E; w_imag[22] = 8'hEF;
w_real[23] = 8'h7E; w_imag[23] = 8'hEE;
w_real[24] = 8'h7E; w_imag[24] = 8'hEE;
w_real[25] = 8'h7E; w_imag[25] = 8'hED;
w_real[26] = 8'h7E; w_imag[26] = 8'hEC;
w_real[27] = 8'h7E; w_imag[27] = 8'hEB;
w_real[28] = 8'h7E; w_imag[28] = 8'hEB;
w_real[29] = 8'h7D; w_imag[29] = 8'hEA;
w_real[30] = 8'h7D; w_imag[30] = 8'hE9;
w_real[31] = 8'h7D; w_imag[31] = 8'hE8;
w_real[32] = 8'h7D; w_imag[32] = 8'hE8;
w_real[33] = 8'h7D; w_imag[33] = 8'hE7;
w_real[34] = 8'h7D; w_imag[34] = 8'hE6;
w_real[35] = 8'h7D; w_imag[35] = 8'hE5;
w_real[36] = 8'h7C; w_imag[36] = 8'hE4;
w_real[37] = 8'h7C; w_imag[37] = 8'hE4;
w_real[38] = 8'h7C; w_imag[38] = 8'hE3;
w_real[39] = 8'h7C; w_imag[39] = 8'hE2;
w_real[40] = 8'h7C; w_imag[40] = 8'hE1;
w_real[41] = 8'h7B; w_imag[41] = 8'hE1;
w_real[42] = 8'h7B; w_imag[42] = 8'hE0;
w_real[43] = 8'h7B; w_imag[43] = 8'hDF;
w_real[44] = 8'h7B; w_imag[44] = 8'hDE;
w_real[45] = 8'h7B; w_imag[45] = 8'hDE;
w_real[46] = 8'h7A; w_imag[46] = 8'hDD;
w_real[47] = 8'h7A; w_imag[47] = 8'hDC;
w_real[48] = 8'h7A; w_imag[48] = 8'hDB;
w_real[49] = 8'h7A; w_imag[49] = 8'hDB;
w_real[50] = 8'h7A; w_imag[50] = 8'hDA;
w_real[51] = 8'h79; w_imag[51] = 8'hD9;
w_real[52] = 8'h79; w_imag[52] = 8'hD8;
w_real[53] = 8'h79; w_imag[53] = 8'hD8;
w_real[54] = 8'h79; w_imag[54] = 8'hD7;
w_real[55] = 8'h78; w_imag[55] = 8'hD6;
w_real[56] = 8'h78; w_imag[56] = 8'hD5;
w_real[57] = 8'h78; w_imag[57] = 8'hD5;
w_real[58] = 8'h77; w_imag[58] = 8'hD4;
w_real[59] = 8'h77; w_imag[59] = 8'hD3;
w_real[60] = 8'h77; w_imag[60] = 8'hD2;
w_real[61] = 8'h77; w_imag[61] = 8'hD2;
w_real[62] = 8'h76; w_imag[62] = 8'hD1;
w_real[63] = 8'h76; w_imag[63] = 8'hD0;
w_real[64] = 8'h76; w_imag[64] = 8'hD0;
w_real[65] = 8'h75; w_imag[65] = 8'hCF;
w_real[66] = 8'h75; w_imag[66] = 8'hCE;
w_real[67] = 8'h75; w_imag[67] = 8'hCD;
w_real[68] = 8'h75; w_imag[68] = 8'hCD;
w_real[69] = 8'h74; w_imag[69] = 8'hCC;
w_real[70] = 8'h74; w_imag[70] = 8'hCB;
w_real[71] = 8'h74; w_imag[71] = 8'hCA;
w_real[72] = 8'h73; w_imag[72] = 8'hCA;
w_real[73] = 8'h73; w_imag[73] = 8'hC9;
w_real[74] = 8'h73; w_imag[74] = 8'hC8;
w_real[75] = 8'h72; w_imag[75] = 8'hC8;
w_real[76] = 8'h72; w_imag[76] = 8'hC7;
w_real[77] = 8'h71; w_imag[77] = 8'hC6;
w_real[78] = 8'h71; w_imag[78] = 8'hC6;
w_real[79] = 8'h71; w_imag[79] = 8'hC5;
w_real[80] = 8'h70; w_imag[80] = 8'hC4;
w_real[81] = 8'h70; w_imag[81] = 8'hC3;
w_real[82] = 8'h70; w_imag[82] = 8'hC3;
w_real[83] = 8'h6F; w_imag[83] = 8'hC2;
w_real[84] = 8'h6F; w_imag[84] = 8'hC1;
w_real[85] = 8'h6E; w_imag[85] = 8'hC1;
w_real[86] = 8'h6E; w_imag[86] = 8'hC0;
w_real[87] = 8'h6E; w_imag[87] = 8'hBF;
w_real[88] = 8'h6D; w_imag[88] = 8'hBF;
w_real[89] = 8'h6D; w_imag[89] = 8'hBE;
w_real[90] = 8'h6C; w_imag[90] = 8'hBD;
w_real[91] = 8'h6C; w_imag[91] = 8'hBD;
w_real[92] = 8'h6C; w_imag[92] = 8'hBC;
w_real[93] = 8'h6B; w_imag[93] = 8'hBB;
w_real[94] = 8'h6B; w_imag[94] = 8'hBB;
w_real[95] = 8'h6A; w_imag[95] = 8'hBA;
w_real[96] = 8'h6A; w_imag[96] = 8'hB9;
w_real[97] = 8'h69; w_imag[97] = 8'hB9;
w_real[98] = 8'h69; w_imag[98] = 8'hB8;
w_real[99] = 8'h69; w_imag[99] = 8'hB7;
w_real[100] = 8'h68; w_imag[100] = 8'hB7;
w_real[101] = 8'h68; w_imag[101] = 8'hB6;
w_real[102] = 8'h67; w_imag[102] = 8'hB6;
w_real[103] = 8'h67; w_imag[103] = 8'hB5;
w_real[104] = 8'h66; w_imag[104] = 8'hB4;
w_real[105] = 8'h66; w_imag[105] = 8'hB4;
w_real[106] = 8'h65; w_imag[106] = 8'hB3;
w_real[107] = 8'h65; w_imag[107] = 8'hB2;
w_real[108] = 8'h64; w_imag[108] = 8'hB2;
w_real[109] = 8'h64; w_imag[109] = 8'hB1;
w_real[110] = 8'h63; w_imag[110] = 8'hB1;
w_real[111] = 8'h63; w_imag[111] = 8'hB0;
w_real[112] = 8'h62; w_imag[112] = 8'hAF;
w_real[113] = 8'h62; w_imag[113] = 8'hAF;
w_real[114] = 8'h61; w_imag[114] = 8'hAE;
w_real[115] = 8'h61; w_imag[115] = 8'hAD;
w_real[116] = 8'h60; w_imag[116] = 8'hAD;
w_real[117] = 8'h60; w_imag[117] = 8'hAC;
w_real[118] = 8'h5F; w_imag[118] = 8'hAC;
w_real[119] = 8'h5F; w_imag[119] = 8'hAB;
w_real[120] = 8'h5E; w_imag[120] = 8'hAB;
w_real[121] = 8'h5E; w_imag[121] = 8'hAA;
w_real[122] = 8'h5D; w_imag[122] = 8'hA9;
w_real[123] = 8'h5D; w_imag[123] = 8'hA9;
w_real[124] = 8'h5C; w_imag[124] = 8'hA8;
w_real[125] = 8'h5C; w_imag[125] = 8'hA8;
w_real[126] = 8'h5B; w_imag[126] = 8'hA7;
w_real[127] = 8'h5B; w_imag[127] = 8'hA7;
w_real[128] = 8'h5A; w_imag[128] = 8'hA6;
w_real[129] = 8'h59; w_imag[129] = 8'hA5;
w_real[130] = 8'h59; w_imag[130] = 8'hA5;
w_real[131] = 8'h58; w_imag[131] = 8'hA4;
w_real[132] = 8'h58; w_imag[132] = 8'hA4;
w_real[133] = 8'h57; w_imag[133] = 8'hA3;
w_real[134] = 8'h57; w_imag[134] = 8'hA3;
w_real[135] = 8'h56; w_imag[135] = 8'hA2;
w_real[136] = 8'h55; w_imag[136] = 8'hA2;
w_real[137] = 8'h55; w_imag[137] = 8'hA1;
w_real[138] = 8'h54; w_imag[138] = 8'hA1;
w_real[139] = 8'h54; w_imag[139] = 8'hA0;
w_real[140] = 8'h53; w_imag[140] = 8'hA0;
w_real[141] = 8'h53; w_imag[141] = 8'h9F;
w_real[142] = 8'h52; w_imag[142] = 8'h9F;
w_real[143] = 8'h51; w_imag[143] = 8'h9E;
w_real[144] = 8'h51; w_imag[144] = 8'h9E;
w_real[145] = 8'h50; w_imag[145] = 8'h9D;
w_real[146] = 8'h4F; w_imag[146] = 8'h9D;
w_real[147] = 8'h4F; w_imag[147] = 8'h9C;
w_real[148] = 8'h4E; w_imag[148] = 8'h9C;
w_real[149] = 8'h4E; w_imag[149] = 8'h9B;
w_real[150] = 8'h4D; w_imag[150] = 8'h9B;
w_real[151] = 8'h4C; w_imag[151] = 8'h9A;
w_real[152] = 8'h4C; w_imag[152] = 8'h9A;
w_real[153] = 8'h4B; w_imag[153] = 8'h99;
w_real[154] = 8'h4A; w_imag[154] = 8'h99;
w_real[155] = 8'h4A; w_imag[155] = 8'h98;
w_real[156] = 8'h49; w_imag[156] = 8'h98;
w_real[157] = 8'h49; w_imag[157] = 8'h97;
w_real[158] = 8'h48; w_imag[158] = 8'h97;
w_real[159] = 8'h47; w_imag[159] = 8'h97;
w_real[160] = 8'h47; w_imag[160] = 8'h96;
w_real[161] = 8'h46; w_imag[161] = 8'h96;
w_real[162] = 8'h45; w_imag[162] = 8'h95;
w_real[163] = 8'h45; w_imag[163] = 8'h95;
w_real[164] = 8'h44; w_imag[164] = 8'h94;
w_real[165] = 8'h43; w_imag[165] = 8'h94;
w_real[166] = 8'h43; w_imag[166] = 8'h94;
w_real[167] = 8'h42; w_imag[167] = 8'h93;
w_real[168] = 8'h41; w_imag[168] = 8'h93;
w_real[169] = 8'h41; w_imag[169] = 8'h92;
w_real[170] = 8'h40; w_imag[170] = 8'h92;
w_real[171] = 8'h3F; w_imag[171] = 8'h92;
w_real[172] = 8'h3F; w_imag[172] = 8'h91;
w_real[173] = 8'h3E; w_imag[173] = 8'h91;
w_real[174] = 8'h3D; w_imag[174] = 8'h90;
w_real[175] = 8'h3D; w_imag[175] = 8'h90;
w_real[176] = 8'h3C; w_imag[176] = 8'h90;
w_real[177] = 8'h3B; w_imag[177] = 8'h8F;
w_real[178] = 8'h3A; w_imag[178] = 8'h8F;
w_real[179] = 8'h3A; w_imag[179] = 8'h8F;
w_real[180] = 8'h39; w_imag[180] = 8'h8E;
w_real[181] = 8'h38; w_imag[181] = 8'h8E;
w_real[182] = 8'h38; w_imag[182] = 8'h8D;
w_real[183] = 8'h37; w_imag[183] = 8'h8D;
w_real[184] = 8'h36; w_imag[184] = 8'h8D;
w_real[185] = 8'h36; w_imag[185] = 8'h8C;
w_real[186] = 8'h35; w_imag[186] = 8'h8C;
w_real[187] = 8'h34; w_imag[187] = 8'h8C;
w_real[188] = 8'h33; w_imag[188] = 8'h8B;
w_real[189] = 8'h33; w_imag[189] = 8'h8B;
w_real[190] = 8'h32; w_imag[190] = 8'h8B;
w_real[191] = 8'h31; w_imag[191] = 8'h8B;
w_real[192] = 8'h30; w_imag[192] = 8'h8A;
w_real[193] = 8'h30; w_imag[193] = 8'h8A;
w_real[194] = 8'h2F; w_imag[194] = 8'h8A;
w_real[195] = 8'h2E; w_imag[195] = 8'h89;
w_real[196] = 8'h2E; w_imag[196] = 8'h89;
w_real[197] = 8'h2D; w_imag[197] = 8'h89;
w_real[198] = 8'h2C; w_imag[198] = 8'h89;
w_real[199] = 8'h2B; w_imag[199] = 8'h88;
w_real[200] = 8'h2B; w_imag[200] = 8'h88;
w_real[201] = 8'h2A; w_imag[201] = 8'h88;
w_real[202] = 8'h29; w_imag[202] = 8'h87;
w_real[203] = 8'h28; w_imag[203] = 8'h87;
w_real[204] = 8'h28; w_imag[204] = 8'h87;
w_real[205] = 8'h27; w_imag[205] = 8'h87;
w_real[206] = 8'h26; w_imag[206] = 8'h86;
w_real[207] = 8'h25; w_imag[207] = 8'h86;
w_real[208] = 8'h25; w_imag[208] = 8'h86;
w_real[209] = 8'h24; w_imag[209] = 8'h86;
w_real[210] = 8'h23; w_imag[210] = 8'h86;
w_real[211] = 8'h22; w_imag[211] = 8'h85;
w_real[212] = 8'h22; w_imag[212] = 8'h85;
w_real[213] = 8'h21; w_imag[213] = 8'h85;
w_real[214] = 8'h20; w_imag[214] = 8'h85;
w_real[215] = 8'h1F; w_imag[215] = 8'h85;
w_real[216] = 8'h1F; w_imag[216] = 8'h84;
w_real[217] = 8'h1E; w_imag[217] = 8'h84;
w_real[218] = 8'h1D; w_imag[218] = 8'h84;
w_real[219] = 8'h1C; w_imag[219] = 8'h84;
w_real[220] = 8'h1C; w_imag[220] = 8'h84;
w_real[221] = 8'h1B; w_imag[221] = 8'h83;
w_real[222] = 8'h1A; w_imag[222] = 8'h83;
w_real[223] = 8'h19; w_imag[223] = 8'h83;
w_real[224] = 8'h18; w_imag[224] = 8'h83;
w_real[225] = 8'h18; w_imag[225] = 8'h83;
w_real[226] = 8'h17; w_imag[226] = 8'h83;
w_real[227] = 8'h16; w_imag[227] = 8'h83;
w_real[228] = 8'h15; w_imag[228] = 8'h82;
w_real[229] = 8'h15; w_imag[229] = 8'h82;
w_real[230] = 8'h14; w_imag[230] = 8'h82;
w_real[231] = 8'h13; w_imag[231] = 8'h82;
w_real[232] = 8'h12; w_imag[232] = 8'h82;
w_real[233] = 8'h12; w_imag[233] = 8'h82;
w_real[234] = 8'h11; w_imag[234] = 8'h82;
w_real[235] = 8'h10; w_imag[235] = 8'h82;
w_real[236] = 8'h0F; w_imag[236] = 8'h81;
w_real[237] = 8'h0E; w_imag[237] = 8'h81;
w_real[238] = 8'h0E; w_imag[238] = 8'h81;
w_real[239] = 8'h0D; w_imag[239] = 8'h81;
w_real[240] = 8'h0C; w_imag[240] = 8'h81;
w_real[241] = 8'h0B; w_imag[241] = 8'h81;
w_real[242] = 8'h0A; w_imag[242] = 8'h81;
w_real[243] = 8'h0A; w_imag[243] = 8'h81;
w_real[244] = 8'h09; w_imag[244] = 8'h81;
w_real[245] = 8'h08; w_imag[245] = 8'h81;
w_real[246] = 8'h07; w_imag[246] = 8'h81;
w_real[247] = 8'h07; w_imag[247] = 8'h81;
w_real[248] = 8'h06; w_imag[248] = 8'h81;
w_real[249] = 8'h05; w_imag[249] = 8'h81;
w_real[250] = 8'h04; w_imag[250] = 8'h81;
w_real[251] = 8'h03; w_imag[251] = 8'h81;
w_real[252] = 8'h03; w_imag[252] = 8'h81;
w_real[253] = 8'h02; w_imag[253] = 8'h81;
w_real[254] = 8'h01; w_imag[254] = 8'h81;
w_real[255] = 8'h00; w_imag[255] = 8'h81;
w_real[256] = 8'h00; w_imag[256] = 8'h80;
w_real[257] = 8'h00; w_imag[257] = 8'h81;
w_real[258] = 8'hFF; w_imag[258] = 8'h81;
w_real[259] = 8'hFE; w_imag[259] = 8'h81;
w_real[260] = 8'hFD; w_imag[260] = 8'h81;
w_real[261] = 8'hFD; w_imag[261] = 8'h81;
w_real[262] = 8'hFC; w_imag[262] = 8'h81;
w_real[263] = 8'hFB; w_imag[263] = 8'h81;
w_real[264] = 8'hFA; w_imag[264] = 8'h81;
w_real[265] = 8'hF9; w_imag[265] = 8'h81;
w_real[266] = 8'hF9; w_imag[266] = 8'h81;
w_real[267] = 8'hF8; w_imag[267] = 8'h81;
w_real[268] = 8'hF7; w_imag[268] = 8'h81;
w_real[269] = 8'hF6; w_imag[269] = 8'h81;
w_real[270] = 8'hF6; w_imag[270] = 8'h81;
w_real[271] = 8'hF5; w_imag[271] = 8'h81;
w_real[272] = 8'hF4; w_imag[272] = 8'h81;
w_real[273] = 8'hF3; w_imag[273] = 8'h81;
w_real[274] = 8'hF2; w_imag[274] = 8'h81;
w_real[275] = 8'hF2; w_imag[275] = 8'h81;
w_real[276] = 8'hF1; w_imag[276] = 8'h81;
w_real[277] = 8'hF0; w_imag[277] = 8'h82;
w_real[278] = 8'hEF; w_imag[278] = 8'h82;
w_real[279] = 8'hEE; w_imag[279] = 8'h82;
w_real[280] = 8'hEE; w_imag[280] = 8'h82;
w_real[281] = 8'hED; w_imag[281] = 8'h82;
w_real[282] = 8'hEC; w_imag[282] = 8'h82;
w_real[283] = 8'hEB; w_imag[283] = 8'h82;
w_real[284] = 8'hEB; w_imag[284] = 8'h82;
w_real[285] = 8'hEA; w_imag[285] = 8'h83;
w_real[286] = 8'hE9; w_imag[286] = 8'h83;
w_real[287] = 8'hE8; w_imag[287] = 8'h83;
w_real[288] = 8'hE8; w_imag[288] = 8'h83;
w_real[289] = 8'hE7; w_imag[289] = 8'h83;
w_real[290] = 8'hE6; w_imag[290] = 8'h83;
w_real[291] = 8'hE5; w_imag[291] = 8'h83;
w_real[292] = 8'hE4; w_imag[292] = 8'h84;
w_real[293] = 8'hE4; w_imag[293] = 8'h84;
w_real[294] = 8'hE3; w_imag[294] = 8'h84;
w_real[295] = 8'hE2; w_imag[295] = 8'h84;
w_real[296] = 8'hE1; w_imag[296] = 8'h84;
w_real[297] = 8'hE1; w_imag[297] = 8'h85;
w_real[298] = 8'hE0; w_imag[298] = 8'h85;
w_real[299] = 8'hDF; w_imag[299] = 8'h85;
w_real[300] = 8'hDE; w_imag[300] = 8'h85;
w_real[301] = 8'hDE; w_imag[301] = 8'h85;
w_real[302] = 8'hDD; w_imag[302] = 8'h86;
w_real[303] = 8'hDC; w_imag[303] = 8'h86;
w_real[304] = 8'hDB; w_imag[304] = 8'h86;
w_real[305] = 8'hDB; w_imag[305] = 8'h86;
w_real[306] = 8'hDA; w_imag[306] = 8'h86;
w_real[307] = 8'hD9; w_imag[307] = 8'h87;
w_real[308] = 8'hD8; w_imag[308] = 8'h87;
w_real[309] = 8'hD8; w_imag[309] = 8'h87;
w_real[310] = 8'hD7; w_imag[310] = 8'h87;
w_real[311] = 8'hD6; w_imag[311] = 8'h88;
w_real[312] = 8'hD5; w_imag[312] = 8'h88;
w_real[313] = 8'hD5; w_imag[313] = 8'h88;
w_real[314] = 8'hD4; w_imag[314] = 8'h89;
w_real[315] = 8'hD3; w_imag[315] = 8'h89;
w_real[316] = 8'hD2; w_imag[316] = 8'h89;
w_real[317] = 8'hD2; w_imag[317] = 8'h89;
w_real[318] = 8'hD1; w_imag[318] = 8'h8A;
w_real[319] = 8'hD0; w_imag[319] = 8'h8A;
w_real[320] = 8'hD0; w_imag[320] = 8'h8A;
w_real[321] = 8'hCF; w_imag[321] = 8'h8B;
w_real[322] = 8'hCE; w_imag[322] = 8'h8B;
w_real[323] = 8'hCD; w_imag[323] = 8'h8B;
w_real[324] = 8'hCD; w_imag[324] = 8'h8B;
w_real[325] = 8'hCC; w_imag[325] = 8'h8C;
w_real[326] = 8'hCB; w_imag[326] = 8'h8C;
w_real[327] = 8'hCA; w_imag[327] = 8'h8C;
w_real[328] = 8'hCA; w_imag[328] = 8'h8D;
w_real[329] = 8'hC9; w_imag[329] = 8'h8D;
w_real[330] = 8'hC8; w_imag[330] = 8'h8D;
w_real[331] = 8'hC8; w_imag[331] = 8'h8E;
w_real[332] = 8'hC7; w_imag[332] = 8'h8E;
w_real[333] = 8'hC6; w_imag[333] = 8'h8F;
w_real[334] = 8'hC6; w_imag[334] = 8'h8F;
w_real[335] = 8'hC5; w_imag[335] = 8'h8F;
w_real[336] = 8'hC4; w_imag[336] = 8'h90;
w_real[337] = 8'hC3; w_imag[337] = 8'h90;
w_real[338] = 8'hC3; w_imag[338] = 8'h90;
w_real[339] = 8'hC2; w_imag[339] = 8'h91;
w_real[340] = 8'hC1; w_imag[340] = 8'h91;
w_real[341] = 8'hC1; w_imag[341] = 8'h92;
w_real[342] = 8'hC0; w_imag[342] = 8'h92;
w_real[343] = 8'hBF; w_imag[343] = 8'h92;
w_real[344] = 8'hBF; w_imag[344] = 8'h93;
w_real[345] = 8'hBE; w_imag[345] = 8'h93;
w_real[346] = 8'hBD; w_imag[346] = 8'h94;
w_real[347] = 8'hBD; w_imag[347] = 8'h94;
w_real[348] = 8'hBC; w_imag[348] = 8'h94;
w_real[349] = 8'hBB; w_imag[349] = 8'h95;
w_real[350] = 8'hBB; w_imag[350] = 8'h95;
w_real[351] = 8'hBA; w_imag[351] = 8'h96;
w_real[352] = 8'hB9; w_imag[352] = 8'h96;
w_real[353] = 8'hB9; w_imag[353] = 8'h97;
w_real[354] = 8'hB8; w_imag[354] = 8'h97;
w_real[355] = 8'hB7; w_imag[355] = 8'h97;
w_real[356] = 8'hB7; w_imag[356] = 8'h98;
w_real[357] = 8'hB6; w_imag[357] = 8'h98;
w_real[358] = 8'hB6; w_imag[358] = 8'h99;
w_real[359] = 8'hB5; w_imag[359] = 8'h99;
w_real[360] = 8'hB4; w_imag[360] = 8'h9A;
w_real[361] = 8'hB4; w_imag[361] = 8'h9A;
w_real[362] = 8'hB3; w_imag[362] = 8'h9B;
w_real[363] = 8'hB2; w_imag[363] = 8'h9B;
w_real[364] = 8'hB2; w_imag[364] = 8'h9C;
w_real[365] = 8'hB1; w_imag[365] = 8'h9C;
w_real[366] = 8'hB1; w_imag[366] = 8'h9D;
w_real[367] = 8'hB0; w_imag[367] = 8'h9D;
w_real[368] = 8'hAF; w_imag[368] = 8'h9E;
w_real[369] = 8'hAF; w_imag[369] = 8'h9E;
w_real[370] = 8'hAE; w_imag[370] = 8'h9F;
w_real[371] = 8'hAD; w_imag[371] = 8'h9F;
w_real[372] = 8'hAD; w_imag[372] = 8'hA0;
w_real[373] = 8'hAC; w_imag[373] = 8'hA0;
w_real[374] = 8'hAC; w_imag[374] = 8'hA1;
w_real[375] = 8'hAB; w_imag[375] = 8'hA1;
w_real[376] = 8'hAB; w_imag[376] = 8'hA2;
w_real[377] = 8'hAA; w_imag[377] = 8'hA2;
w_real[378] = 8'hA9; w_imag[378] = 8'hA3;
w_real[379] = 8'hA9; w_imag[379] = 8'hA3;
w_real[380] = 8'hA8; w_imag[380] = 8'hA4;
w_real[381] = 8'hA8; w_imag[381] = 8'hA4;
w_real[382] = 8'hA7; w_imag[382] = 8'hA5;
w_real[383] = 8'hA7; w_imag[383] = 8'hA5;
w_real[384] = 8'hA6; w_imag[384] = 8'hA6;
w_real[385] = 8'hA5; w_imag[385] = 8'hA7;
w_real[386] = 8'hA5; w_imag[386] = 8'hA7;
w_real[387] = 8'hA4; w_imag[387] = 8'hA8;
w_real[388] = 8'hA4; w_imag[388] = 8'hA8;
w_real[389] = 8'hA3; w_imag[389] = 8'hA9;
w_real[390] = 8'hA3; w_imag[390] = 8'hA9;
w_real[391] = 8'hA2; w_imag[391] = 8'hAA;
w_real[392] = 8'hA2; w_imag[392] = 8'hAB;
w_real[393] = 8'hA1; w_imag[393] = 8'hAB;
w_real[394] = 8'hA1; w_imag[394] = 8'hAC;
w_real[395] = 8'hA0; w_imag[395] = 8'hAC;
w_real[396] = 8'hA0; w_imag[396] = 8'hAD;
w_real[397] = 8'h9F; w_imag[397] = 8'hAD;
w_real[398] = 8'h9F; w_imag[398] = 8'hAE;
w_real[399] = 8'h9E; w_imag[399] = 8'hAF;
w_real[400] = 8'h9E; w_imag[400] = 8'hAF;
w_real[401] = 8'h9D; w_imag[401] = 8'hB0;
w_real[402] = 8'h9D; w_imag[402] = 8'hB1;
w_real[403] = 8'h9C; w_imag[403] = 8'hB1;
w_real[404] = 8'h9C; w_imag[404] = 8'hB2;
w_real[405] = 8'h9B; w_imag[405] = 8'hB2;
w_real[406] = 8'h9B; w_imag[406] = 8'hB3;
w_real[407] = 8'h9A; w_imag[407] = 8'hB4;
w_real[408] = 8'h9A; w_imag[408] = 8'hB4;
w_real[409] = 8'h99; w_imag[409] = 8'hB5;
w_real[410] = 8'h99; w_imag[410] = 8'hB6;
w_real[411] = 8'h98; w_imag[411] = 8'hB6;
w_real[412] = 8'h98; w_imag[412] = 8'hB7;
w_real[413] = 8'h97; w_imag[413] = 8'hB7;
w_real[414] = 8'h97; w_imag[414] = 8'hB8;
w_real[415] = 8'h97; w_imag[415] = 8'hB9;
w_real[416] = 8'h96; w_imag[416] = 8'hB9;
w_real[417] = 8'h96; w_imag[417] = 8'hBA;
w_real[418] = 8'h95; w_imag[418] = 8'hBB;
w_real[419] = 8'h95; w_imag[419] = 8'hBB;
w_real[420] = 8'h94; w_imag[420] = 8'hBC;
w_real[421] = 8'h94; w_imag[421] = 8'hBD;
w_real[422] = 8'h94; w_imag[422] = 8'hBD;
w_real[423] = 8'h93; w_imag[423] = 8'hBE;
w_real[424] = 8'h93; w_imag[424] = 8'hBF;
w_real[425] = 8'h92; w_imag[425] = 8'hBF;
w_real[426] = 8'h92; w_imag[426] = 8'hC0;
w_real[427] = 8'h92; w_imag[427] = 8'hC1;
w_real[428] = 8'h91; w_imag[428] = 8'hC1;
w_real[429] = 8'h91; w_imag[429] = 8'hC2;
w_real[430] = 8'h90; w_imag[430] = 8'hC3;
w_real[431] = 8'h90; w_imag[431] = 8'hC3;
w_real[432] = 8'h90; w_imag[432] = 8'hC4;
w_real[433] = 8'h8F; w_imag[433] = 8'hC5;
w_real[434] = 8'h8F; w_imag[434] = 8'hC6;
w_real[435] = 8'h8F; w_imag[435] = 8'hC6;
w_real[436] = 8'h8E; w_imag[436] = 8'hC7;
w_real[437] = 8'h8E; w_imag[437] = 8'hC8;
w_real[438] = 8'h8D; w_imag[438] = 8'hC8;
w_real[439] = 8'h8D; w_imag[439] = 8'hC9;
w_real[440] = 8'h8D; w_imag[440] = 8'hCA;
w_real[441] = 8'h8C; w_imag[441] = 8'hCA;
w_real[442] = 8'h8C; w_imag[442] = 8'hCB;
w_real[443] = 8'h8C; w_imag[443] = 8'hCC;
w_real[444] = 8'h8B; w_imag[444] = 8'hCD;
w_real[445] = 8'h8B; w_imag[445] = 8'hCD;
w_real[446] = 8'h8B; w_imag[446] = 8'hCE;
w_real[447] = 8'h8B; w_imag[447] = 8'hCF;
w_real[448] = 8'h8A; w_imag[448] = 8'hD0;
w_real[449] = 8'h8A; w_imag[449] = 8'hD0;
w_real[450] = 8'h8A; w_imag[450] = 8'hD1;
w_real[451] = 8'h89; w_imag[451] = 8'hD2;
w_real[452] = 8'h89; w_imag[452] = 8'hD2;
w_real[453] = 8'h89; w_imag[453] = 8'hD3;
w_real[454] = 8'h89; w_imag[454] = 8'hD4;
w_real[455] = 8'h88; w_imag[455] = 8'hD5;
w_real[456] = 8'h88; w_imag[456] = 8'hD5;
w_real[457] = 8'h88; w_imag[457] = 8'hD6;
w_real[458] = 8'h87; w_imag[458] = 8'hD7;
w_real[459] = 8'h87; w_imag[459] = 8'hD8;
w_real[460] = 8'h87; w_imag[460] = 8'hD8;
w_real[461] = 8'h87; w_imag[461] = 8'hD9;
w_real[462] = 8'h86; w_imag[462] = 8'hDA;
w_real[463] = 8'h86; w_imag[463] = 8'hDB;
w_real[464] = 8'h86; w_imag[464] = 8'hDB;
w_real[465] = 8'h86; w_imag[465] = 8'hDC;
w_real[466] = 8'h86; w_imag[466] = 8'hDD;
w_real[467] = 8'h85; w_imag[467] = 8'hDE;
w_real[468] = 8'h85; w_imag[468] = 8'hDE;
w_real[469] = 8'h85; w_imag[469] = 8'hDF;
w_real[470] = 8'h85; w_imag[470] = 8'hE0;
w_real[471] = 8'h85; w_imag[471] = 8'hE1;
w_real[472] = 8'h84; w_imag[472] = 8'hE1;
w_real[473] = 8'h84; w_imag[473] = 8'hE2;
w_real[474] = 8'h84; w_imag[474] = 8'hE3;
w_real[475] = 8'h84; w_imag[475] = 8'hE4;
w_real[476] = 8'h84; w_imag[476] = 8'hE4;
w_real[477] = 8'h83; w_imag[477] = 8'hE5;
w_real[478] = 8'h83; w_imag[478] = 8'hE6;
w_real[479] = 8'h83; w_imag[479] = 8'hE7;
w_real[480] = 8'h83; w_imag[480] = 8'hE8;
w_real[481] = 8'h83; w_imag[481] = 8'hE8;
w_real[482] = 8'h83; w_imag[482] = 8'hE9;
w_real[483] = 8'h83; w_imag[483] = 8'hEA;
w_real[484] = 8'h82; w_imag[484] = 8'hEB;
w_real[485] = 8'h82; w_imag[485] = 8'hEB;
w_real[486] = 8'h82; w_imag[486] = 8'hEC;
w_real[487] = 8'h82; w_imag[487] = 8'hED;
w_real[488] = 8'h82; w_imag[488] = 8'hEE;
w_real[489] = 8'h82; w_imag[489] = 8'hEE;
w_real[490] = 8'h82; w_imag[490] = 8'hEF;
w_real[491] = 8'h82; w_imag[491] = 8'hF0;
w_real[492] = 8'h81; w_imag[492] = 8'hF1;
w_real[493] = 8'h81; w_imag[493] = 8'hF2;
w_real[494] = 8'h81; w_imag[494] = 8'hF2;
w_real[495] = 8'h81; w_imag[495] = 8'hF3;
w_real[496] = 8'h81; w_imag[496] = 8'hF4;
w_real[497] = 8'h81; w_imag[497] = 8'hF5;
w_real[498] = 8'h81; w_imag[498] = 8'hF6;
w_real[499] = 8'h81; w_imag[499] = 8'hF6;
w_real[500] = 8'h81; w_imag[500] = 8'hF7;
w_real[501] = 8'h81; w_imag[501] = 8'hF8;
w_real[502] = 8'h81; w_imag[502] = 8'hF9;
w_real[503] = 8'h81; w_imag[503] = 8'hF9;
w_real[504] = 8'h81; w_imag[504] = 8'hFA;
w_real[505] = 8'h81; w_imag[505] = 8'hFB;
w_real[506] = 8'h81; w_imag[506] = 8'hFC;
w_real[507] = 8'h81; w_imag[507] = 8'hFD;
w_real[508] = 8'h81; w_imag[508] = 8'hFD;
w_real[509] = 8'h81; w_imag[509] = 8'hFE;
w_real[510] = 8'h81; w_imag[510] = 8'hFF;
w_real[511] = 8'h81; w_imag[511] = 8'h00;
w_real[512] = 8'h80; w_imag[512] = 8'h00;
w_real[513] = 8'h81; w_imag[513] = 8'h00;
w_real[514] = 8'h81; w_imag[514] = 8'h01;
w_real[515] = 8'h81; w_imag[515] = 8'h02;
w_real[516] = 8'h81; w_imag[516] = 8'h03;
w_real[517] = 8'h81; w_imag[517] = 8'h03;
w_real[518] = 8'h81; w_imag[518] = 8'h04;
w_real[519] = 8'h81; w_imag[519] = 8'h05;
w_real[520] = 8'h81; w_imag[520] = 8'h06;
w_real[521] = 8'h81; w_imag[521] = 8'h07;
w_real[522] = 8'h81; w_imag[522] = 8'h07;
w_real[523] = 8'h81; w_imag[523] = 8'h08;
w_real[524] = 8'h81; w_imag[524] = 8'h09;
w_real[525] = 8'h81; w_imag[525] = 8'h0A;
w_real[526] = 8'h81; w_imag[526] = 8'h0A;
w_real[527] = 8'h81; w_imag[527] = 8'h0B;
w_real[528] = 8'h81; w_imag[528] = 8'h0C;
w_real[529] = 8'h81; w_imag[529] = 8'h0D;
w_real[530] = 8'h81; w_imag[530] = 8'h0E;
w_real[531] = 8'h81; w_imag[531] = 8'h0E;
w_real[532] = 8'h81; w_imag[532] = 8'h0F;
w_real[533] = 8'h82; w_imag[533] = 8'h10;
w_real[534] = 8'h82; w_imag[534] = 8'h11;
w_real[535] = 8'h82; w_imag[535] = 8'h12;
w_real[536] = 8'h82; w_imag[536] = 8'h12;
w_real[537] = 8'h82; w_imag[537] = 8'h13;
w_real[538] = 8'h82; w_imag[538] = 8'h14;
w_real[539] = 8'h82; w_imag[539] = 8'h15;
w_real[540] = 8'h82; w_imag[540] = 8'h15;
w_real[541] = 8'h83; w_imag[541] = 8'h16;
w_real[542] = 8'h83; w_imag[542] = 8'h17;
w_real[543] = 8'h83; w_imag[543] = 8'h18;
w_real[544] = 8'h83; w_imag[544] = 8'h18;
w_real[545] = 8'h83; w_imag[545] = 8'h19;
w_real[546] = 8'h83; w_imag[546] = 8'h1A;
w_real[547] = 8'h83; w_imag[547] = 8'h1B;
w_real[548] = 8'h84; w_imag[548] = 8'h1C;
w_real[549] = 8'h84; w_imag[549] = 8'h1C;
w_real[550] = 8'h84; w_imag[550] = 8'h1D;
w_real[551] = 8'h84; w_imag[551] = 8'h1E;
w_real[552] = 8'h84; w_imag[552] = 8'h1F;
w_real[553] = 8'h85; w_imag[553] = 8'h1F;
w_real[554] = 8'h85; w_imag[554] = 8'h20;
w_real[555] = 8'h85; w_imag[555] = 8'h21;
w_real[556] = 8'h85; w_imag[556] = 8'h22;
w_real[557] = 8'h85; w_imag[557] = 8'h22;
w_real[558] = 8'h86; w_imag[558] = 8'h23;
w_real[559] = 8'h86; w_imag[559] = 8'h24;
w_real[560] = 8'h86; w_imag[560] = 8'h25;
w_real[561] = 8'h86; w_imag[561] = 8'h25;
w_real[562] = 8'h86; w_imag[562] = 8'h26;
w_real[563] = 8'h87; w_imag[563] = 8'h27;
w_real[564] = 8'h87; w_imag[564] = 8'h28;
w_real[565] = 8'h87; w_imag[565] = 8'h28;
w_real[566] = 8'h87; w_imag[566] = 8'h29;
w_real[567] = 8'h88; w_imag[567] = 8'h2A;
w_real[568] = 8'h88; w_imag[568] = 8'h2B;
w_real[569] = 8'h88; w_imag[569] = 8'h2B;
w_real[570] = 8'h89; w_imag[570] = 8'h2C;
w_real[571] = 8'h89; w_imag[571] = 8'h2D;
w_real[572] = 8'h89; w_imag[572] = 8'h2E;
w_real[573] = 8'h89; w_imag[573] = 8'h2E;
w_real[574] = 8'h8A; w_imag[574] = 8'h2F;
w_real[575] = 8'h8A; w_imag[575] = 8'h30;
w_real[576] = 8'h8A; w_imag[576] = 8'h30;
w_real[577] = 8'h8B; w_imag[577] = 8'h31;
w_real[578] = 8'h8B; w_imag[578] = 8'h32;
w_real[579] = 8'h8B; w_imag[579] = 8'h33;
w_real[580] = 8'h8B; w_imag[580] = 8'h33;
w_real[581] = 8'h8C; w_imag[581] = 8'h34;
w_real[582] = 8'h8C; w_imag[582] = 8'h35;
w_real[583] = 8'h8C; w_imag[583] = 8'h36;
w_real[584] = 8'h8D; w_imag[584] = 8'h36;
w_real[585] = 8'h8D; w_imag[585] = 8'h37;
w_real[586] = 8'h8D; w_imag[586] = 8'h38;
w_real[587] = 8'h8E; w_imag[587] = 8'h38;
w_real[588] = 8'h8E; w_imag[588] = 8'h39;
w_real[589] = 8'h8F; w_imag[589] = 8'h3A;
w_real[590] = 8'h8F; w_imag[590] = 8'h3A;
w_real[591] = 8'h8F; w_imag[591] = 8'h3B;
w_real[592] = 8'h90; w_imag[592] = 8'h3C;
w_real[593] = 8'h90; w_imag[593] = 8'h3D;
w_real[594] = 8'h90; w_imag[594] = 8'h3D;
w_real[595] = 8'h91; w_imag[595] = 8'h3E;
w_real[596] = 8'h91; w_imag[596] = 8'h3F;
w_real[597] = 8'h92; w_imag[597] = 8'h3F;
w_real[598] = 8'h92; w_imag[598] = 8'h40;
w_real[599] = 8'h92; w_imag[599] = 8'h41;
w_real[600] = 8'h93; w_imag[600] = 8'h41;
w_real[601] = 8'h93; w_imag[601] = 8'h42;
w_real[602] = 8'h94; w_imag[602] = 8'h43;
w_real[603] = 8'h94; w_imag[603] = 8'h43;
w_real[604] = 8'h94; w_imag[604] = 8'h44;
w_real[605] = 8'h95; w_imag[605] = 8'h45;
w_real[606] = 8'h95; w_imag[606] = 8'h45;
w_real[607] = 8'h96; w_imag[607] = 8'h46;
w_real[608] = 8'h96; w_imag[608] = 8'h47;
w_real[609] = 8'h97; w_imag[609] = 8'h47;
w_real[610] = 8'h97; w_imag[610] = 8'h48;
w_real[611] = 8'h97; w_imag[611] = 8'h49;
w_real[612] = 8'h98; w_imag[612] = 8'h49;
w_real[613] = 8'h98; w_imag[613] = 8'h4A;
w_real[614] = 8'h99; w_imag[614] = 8'h4A;
w_real[615] = 8'h99; w_imag[615] = 8'h4B;
w_real[616] = 8'h9A; w_imag[616] = 8'h4C;
w_real[617] = 8'h9A; w_imag[617] = 8'h4C;
w_real[618] = 8'h9B; w_imag[618] = 8'h4D;
w_real[619] = 8'h9B; w_imag[619] = 8'h4E;
w_real[620] = 8'h9C; w_imag[620] = 8'h4E;
w_real[621] = 8'h9C; w_imag[621] = 8'h4F;
w_real[622] = 8'h9D; w_imag[622] = 8'h4F;
w_real[623] = 8'h9D; w_imag[623] = 8'h50;
w_real[624] = 8'h9E; w_imag[624] = 8'h51;
w_real[625] = 8'h9E; w_imag[625] = 8'h51;
w_real[626] = 8'h9F; w_imag[626] = 8'h52;
w_real[627] = 8'h9F; w_imag[627] = 8'h53;
w_real[628] = 8'hA0; w_imag[628] = 8'h53;
w_real[629] = 8'hA0; w_imag[629] = 8'h54;
w_real[630] = 8'hA1; w_imag[630] = 8'h54;
w_real[631] = 8'hA1; w_imag[631] = 8'h55;
w_real[632] = 8'hA2; w_imag[632] = 8'h55;
w_real[633] = 8'hA2; w_imag[633] = 8'h56;
w_real[634] = 8'hA3; w_imag[634] = 8'h57;
w_real[635] = 8'hA3; w_imag[635] = 8'h57;
w_real[636] = 8'hA4; w_imag[636] = 8'h58;
w_real[637] = 8'hA4; w_imag[637] = 8'h58;
w_real[638] = 8'hA5; w_imag[638] = 8'h59;
w_real[639] = 8'hA5; w_imag[639] = 8'h59;
w_real[640] = 8'hA6; w_imag[640] = 8'h5A;
w_real[641] = 8'hA7; w_imag[641] = 8'h5B;
w_real[642] = 8'hA7; w_imag[642] = 8'h5B;
w_real[643] = 8'hA8; w_imag[643] = 8'h5C;
w_real[644] = 8'hA8; w_imag[644] = 8'h5C;
w_real[645] = 8'hA9; w_imag[645] = 8'h5D;
w_real[646] = 8'hA9; w_imag[646] = 8'h5D;
w_real[647] = 8'hAA; w_imag[647] = 8'h5E;
w_real[648] = 8'hAB; w_imag[648] = 8'h5E;
w_real[649] = 8'hAB; w_imag[649] = 8'h5F;
w_real[650] = 8'hAC; w_imag[650] = 8'h5F;
w_real[651] = 8'hAC; w_imag[651] = 8'h60;
w_real[652] = 8'hAD; w_imag[652] = 8'h60;
w_real[653] = 8'hAD; w_imag[653] = 8'h61;
w_real[654] = 8'hAE; w_imag[654] = 8'h61;
w_real[655] = 8'hAF; w_imag[655] = 8'h62;
w_real[656] = 8'hAF; w_imag[656] = 8'h62;
w_real[657] = 8'hB0; w_imag[657] = 8'h63;
w_real[658] = 8'hB1; w_imag[658] = 8'h63;
w_real[659] = 8'hB1; w_imag[659] = 8'h64;
w_real[660] = 8'hB2; w_imag[660] = 8'h64;
w_real[661] = 8'hB2; w_imag[661] = 8'h65;
w_real[662] = 8'hB3; w_imag[662] = 8'h65;
w_real[663] = 8'hB4; w_imag[663] = 8'h66;
w_real[664] = 8'hB4; w_imag[664] = 8'h66;
w_real[665] = 8'hB5; w_imag[665] = 8'h67;
w_real[666] = 8'hB6; w_imag[666] = 8'h67;
w_real[667] = 8'hB6; w_imag[667] = 8'h68;
w_real[668] = 8'hB7; w_imag[668] = 8'h68;
w_real[669] = 8'hB7; w_imag[669] = 8'h69;
w_real[670] = 8'hB8; w_imag[670] = 8'h69;
w_real[671] = 8'hB9; w_imag[671] = 8'h69;
w_real[672] = 8'hB9; w_imag[672] = 8'h6A;
w_real[673] = 8'hBA; w_imag[673] = 8'h6A;
w_real[674] = 8'hBB; w_imag[674] = 8'h6B;
w_real[675] = 8'hBB; w_imag[675] = 8'h6B;
w_real[676] = 8'hBC; w_imag[676] = 8'h6C;
w_real[677] = 8'hBD; w_imag[677] = 8'h6C;
w_real[678] = 8'hBD; w_imag[678] = 8'h6C;
w_real[679] = 8'hBE; w_imag[679] = 8'h6D;
w_real[680] = 8'hBF; w_imag[680] = 8'h6D;
w_real[681] = 8'hBF; w_imag[681] = 8'h6E;
w_real[682] = 8'hC0; w_imag[682] = 8'h6E;
w_real[683] = 8'hC1; w_imag[683] = 8'h6E;
w_real[684] = 8'hC1; w_imag[684] = 8'h6F;
w_real[685] = 8'hC2; w_imag[685] = 8'h6F;
w_real[686] = 8'hC3; w_imag[686] = 8'h70;
w_real[687] = 8'hC3; w_imag[687] = 8'h70;
w_real[688] = 8'hC4; w_imag[688] = 8'h70;
w_real[689] = 8'hC5; w_imag[689] = 8'h71;
w_real[690] = 8'hC6; w_imag[690] = 8'h71;
w_real[691] = 8'hC6; w_imag[691] = 8'h71;
w_real[692] = 8'hC7; w_imag[692] = 8'h72;
w_real[693] = 8'hC8; w_imag[693] = 8'h72;
w_real[694] = 8'hC8; w_imag[694] = 8'h73;
w_real[695] = 8'hC9; w_imag[695] = 8'h73;
w_real[696] = 8'hCA; w_imag[696] = 8'h73;
w_real[697] = 8'hCA; w_imag[697] = 8'h74;
w_real[698] = 8'hCB; w_imag[698] = 8'h74;
w_real[699] = 8'hCC; w_imag[699] = 8'h74;
w_real[700] = 8'hCD; w_imag[700] = 8'h75;
w_real[701] = 8'hCD; w_imag[701] = 8'h75;
w_real[702] = 8'hCE; w_imag[702] = 8'h75;
w_real[703] = 8'hCF; w_imag[703] = 8'h75;
w_real[704] = 8'hD0; w_imag[704] = 8'h76;
w_real[705] = 8'hD0; w_imag[705] = 8'h76;
w_real[706] = 8'hD1; w_imag[706] = 8'h76;
w_real[707] = 8'hD2; w_imag[707] = 8'h77;
w_real[708] = 8'hD2; w_imag[708] = 8'h77;
w_real[709] = 8'hD3; w_imag[709] = 8'h77;
w_real[710] = 8'hD4; w_imag[710] = 8'h77;
w_real[711] = 8'hD5; w_imag[711] = 8'h78;
w_real[712] = 8'hD5; w_imag[712] = 8'h78;
w_real[713] = 8'hD6; w_imag[713] = 8'h78;
w_real[714] = 8'hD7; w_imag[714] = 8'h79;
w_real[715] = 8'hD8; w_imag[715] = 8'h79;
w_real[716] = 8'hD8; w_imag[716] = 8'h79;
w_real[717] = 8'hD9; w_imag[717] = 8'h79;
w_real[718] = 8'hDA; w_imag[718] = 8'h7A;
w_real[719] = 8'hDB; w_imag[719] = 8'h7A;
w_real[720] = 8'hDB; w_imag[720] = 8'h7A;
w_real[721] = 8'hDC; w_imag[721] = 8'h7A;
w_real[722] = 8'hDD; w_imag[722] = 8'h7A;
w_real[723] = 8'hDE; w_imag[723] = 8'h7B;
w_real[724] = 8'hDE; w_imag[724] = 8'h7B;
w_real[725] = 8'hDF; w_imag[725] = 8'h7B;
w_real[726] = 8'hE0; w_imag[726] = 8'h7B;
w_real[727] = 8'hE1; w_imag[727] = 8'h7B;
w_real[728] = 8'hE1; w_imag[728] = 8'h7C;
w_real[729] = 8'hE2; w_imag[729] = 8'h7C;
w_real[730] = 8'hE3; w_imag[730] = 8'h7C;
w_real[731] = 8'hE4; w_imag[731] = 8'h7C;
w_real[732] = 8'hE4; w_imag[732] = 8'h7C;
w_real[733] = 8'hE5; w_imag[733] = 8'h7D;
w_real[734] = 8'hE6; w_imag[734] = 8'h7D;
w_real[735] = 8'hE7; w_imag[735] = 8'h7D;
w_real[736] = 8'hE8; w_imag[736] = 8'h7D;
w_real[737] = 8'hE8; w_imag[737] = 8'h7D;
w_real[738] = 8'hE9; w_imag[738] = 8'h7D;
w_real[739] = 8'hEA; w_imag[739] = 8'h7D;
w_real[740] = 8'hEB; w_imag[740] = 8'h7E;
w_real[741] = 8'hEB; w_imag[741] = 8'h7E;
w_real[742] = 8'hEC; w_imag[742] = 8'h7E;
w_real[743] = 8'hED; w_imag[743] = 8'h7E;
w_real[744] = 8'hEE; w_imag[744] = 8'h7E;
w_real[745] = 8'hEE; w_imag[745] = 8'h7E;
w_real[746] = 8'hEF; w_imag[746] = 8'h7E;
w_real[747] = 8'hF0; w_imag[747] = 8'h7E;
w_real[748] = 8'hF1; w_imag[748] = 8'h7F;
w_real[749] = 8'hF2; w_imag[749] = 8'h7F;
w_real[750] = 8'hF2; w_imag[750] = 8'h7F;
w_real[751] = 8'hF3; w_imag[751] = 8'h7F;
w_real[752] = 8'hF4; w_imag[752] = 8'h7F;
w_real[753] = 8'hF5; w_imag[753] = 8'h7F;
w_real[754] = 8'hF6; w_imag[754] = 8'h7F;
w_real[755] = 8'hF6; w_imag[755] = 8'h7F;
w_real[756] = 8'hF7; w_imag[756] = 8'h7F;
w_real[757] = 8'hF8; w_imag[757] = 8'h7F;
w_real[758] = 8'hF9; w_imag[758] = 8'h7F;
w_real[759] = 8'hF9; w_imag[759] = 8'h7F;
w_real[760] = 8'hFA; w_imag[760] = 8'h7F;
w_real[761] = 8'hFB; w_imag[761] = 8'h7F;
w_real[762] = 8'hFC; w_imag[762] = 8'h7F;
w_real[763] = 8'hFD; w_imag[763] = 8'h7F;
w_real[764] = 8'hFD; w_imag[764] = 8'h7F;
w_real[765] = 8'hFE; w_imag[765] = 8'h7F;
w_real[766] = 8'hFF; w_imag[766] = 8'h7F;
w_real[767] = 8'h00; w_imag[767] = 8'h7F;
w_real[768] = 8'h00; w_imag[768] = 8'h7F;
w_real[769] = 8'h00; w_imag[769] = 8'h7F;
w_real[770] = 8'h01; w_imag[770] = 8'h7F;
w_real[771] = 8'h02; w_imag[771] = 8'h7F;
w_real[772] = 8'h03; w_imag[772] = 8'h7F;
w_real[773] = 8'h03; w_imag[773] = 8'h7F;
w_real[774] = 8'h04; w_imag[774] = 8'h7F;
w_real[775] = 8'h05; w_imag[775] = 8'h7F;
w_real[776] = 8'h06; w_imag[776] = 8'h7F;
w_real[777] = 8'h07; w_imag[777] = 8'h7F;
w_real[778] = 8'h07; w_imag[778] = 8'h7F;
w_real[779] = 8'h08; w_imag[779] = 8'h7F;
w_real[780] = 8'h09; w_imag[780] = 8'h7F;
w_real[781] = 8'h0A; w_imag[781] = 8'h7F;
w_real[782] = 8'h0A; w_imag[782] = 8'h7F;
w_real[783] = 8'h0B; w_imag[783] = 8'h7F;
w_real[784] = 8'h0C; w_imag[784] = 8'h7F;
w_real[785] = 8'h0D; w_imag[785] = 8'h7F;
w_real[786] = 8'h0E; w_imag[786] = 8'h7F;
w_real[787] = 8'h0E; w_imag[787] = 8'h7F;
w_real[788] = 8'h0F; w_imag[788] = 8'h7F;
w_real[789] = 8'h10; w_imag[789] = 8'h7E;
w_real[790] = 8'h11; w_imag[790] = 8'h7E;
w_real[791] = 8'h12; w_imag[791] = 8'h7E;
w_real[792] = 8'h12; w_imag[792] = 8'h7E;
w_real[793] = 8'h13; w_imag[793] = 8'h7E;
w_real[794] = 8'h14; w_imag[794] = 8'h7E;
w_real[795] = 8'h15; w_imag[795] = 8'h7E;
w_real[796] = 8'h15; w_imag[796] = 8'h7E;
w_real[797] = 8'h16; w_imag[797] = 8'h7D;
w_real[798] = 8'h17; w_imag[798] = 8'h7D;
w_real[799] = 8'h18; w_imag[799] = 8'h7D;
w_real[800] = 8'h18; w_imag[800] = 8'h7D;
w_real[801] = 8'h19; w_imag[801] = 8'h7D;
w_real[802] = 8'h1A; w_imag[802] = 8'h7D;
w_real[803] = 8'h1B; w_imag[803] = 8'h7D;
w_real[804] = 8'h1C; w_imag[804] = 8'h7C;
w_real[805] = 8'h1C; w_imag[805] = 8'h7C;
w_real[806] = 8'h1D; w_imag[806] = 8'h7C;
w_real[807] = 8'h1E; w_imag[807] = 8'h7C;
w_real[808] = 8'h1F; w_imag[808] = 8'h7C;
w_real[809] = 8'h1F; w_imag[809] = 8'h7B;
w_real[810] = 8'h20; w_imag[810] = 8'h7B;
w_real[811] = 8'h21; w_imag[811] = 8'h7B;
w_real[812] = 8'h22; w_imag[812] = 8'h7B;
w_real[813] = 8'h22; w_imag[813] = 8'h7B;
w_real[814] = 8'h23; w_imag[814] = 8'h7A;
w_real[815] = 8'h24; w_imag[815] = 8'h7A;
w_real[816] = 8'h25; w_imag[816] = 8'h7A;
w_real[817] = 8'h25; w_imag[817] = 8'h7A;
w_real[818] = 8'h26; w_imag[818] = 8'h7A;
w_real[819] = 8'h27; w_imag[819] = 8'h79;
w_real[820] = 8'h28; w_imag[820] = 8'h79;
w_real[821] = 8'h28; w_imag[821] = 8'h79;
w_real[822] = 8'h29; w_imag[822] = 8'h79;
w_real[823] = 8'h2A; w_imag[823] = 8'h78;
w_real[824] = 8'h2B; w_imag[824] = 8'h78;
w_real[825] = 8'h2B; w_imag[825] = 8'h78;
w_real[826] = 8'h2C; w_imag[826] = 8'h77;
w_real[827] = 8'h2D; w_imag[827] = 8'h77;
w_real[828] = 8'h2E; w_imag[828] = 8'h77;
w_real[829] = 8'h2E; w_imag[829] = 8'h77;
w_real[830] = 8'h2F; w_imag[830] = 8'h76;
w_real[831] = 8'h30; w_imag[831] = 8'h76;
w_real[832] = 8'h30; w_imag[832] = 8'h76;
w_real[833] = 8'h31; w_imag[833] = 8'h75;
w_real[834] = 8'h32; w_imag[834] = 8'h75;
w_real[835] = 8'h33; w_imag[835] = 8'h75;
w_real[836] = 8'h33; w_imag[836] = 8'h75;
w_real[837] = 8'h34; w_imag[837] = 8'h74;
w_real[838] = 8'h35; w_imag[838] = 8'h74;
w_real[839] = 8'h36; w_imag[839] = 8'h74;
w_real[840] = 8'h36; w_imag[840] = 8'h73;
w_real[841] = 8'h37; w_imag[841] = 8'h73;
w_real[842] = 8'h38; w_imag[842] = 8'h73;
w_real[843] = 8'h38; w_imag[843] = 8'h72;
w_real[844] = 8'h39; w_imag[844] = 8'h72;
w_real[845] = 8'h3A; w_imag[845] = 8'h71;
w_real[846] = 8'h3A; w_imag[846] = 8'h71;
w_real[847] = 8'h3B; w_imag[847] = 8'h71;
w_real[848] = 8'h3C; w_imag[848] = 8'h70;
w_real[849] = 8'h3D; w_imag[849] = 8'h70;
w_real[850] = 8'h3D; w_imag[850] = 8'h70;
w_real[851] = 8'h3E; w_imag[851] = 8'h6F;
w_real[852] = 8'h3F; w_imag[852] = 8'h6F;
w_real[853] = 8'h3F; w_imag[853] = 8'h6E;
w_real[854] = 8'h40; w_imag[854] = 8'h6E;
w_real[855] = 8'h41; w_imag[855] = 8'h6E;
w_real[856] = 8'h41; w_imag[856] = 8'h6D;
w_real[857] = 8'h42; w_imag[857] = 8'h6D;
w_real[858] = 8'h43; w_imag[858] = 8'h6C;
w_real[859] = 8'h43; w_imag[859] = 8'h6C;
w_real[860] = 8'h44; w_imag[860] = 8'h6C;
w_real[861] = 8'h45; w_imag[861] = 8'h6B;
w_real[862] = 8'h45; w_imag[862] = 8'h6B;
w_real[863] = 8'h46; w_imag[863] = 8'h6A;
w_real[864] = 8'h47; w_imag[864] = 8'h6A;
w_real[865] = 8'h47; w_imag[865] = 8'h69;
w_real[866] = 8'h48; w_imag[866] = 8'h69;
w_real[867] = 8'h49; w_imag[867] = 8'h69;
w_real[868] = 8'h49; w_imag[868] = 8'h68;
w_real[869] = 8'h4A; w_imag[869] = 8'h68;
w_real[870] = 8'h4A; w_imag[870] = 8'h67;
w_real[871] = 8'h4B; w_imag[871] = 8'h67;
w_real[872] = 8'h4C; w_imag[872] = 8'h66;
w_real[873] = 8'h4C; w_imag[873] = 8'h66;
w_real[874] = 8'h4D; w_imag[874] = 8'h65;
w_real[875] = 8'h4E; w_imag[875] = 8'h65;
w_real[876] = 8'h4E; w_imag[876] = 8'h64;
w_real[877] = 8'h4F; w_imag[877] = 8'h64;
w_real[878] = 8'h4F; w_imag[878] = 8'h63;
w_real[879] = 8'h50; w_imag[879] = 8'h63;
w_real[880] = 8'h51; w_imag[880] = 8'h62;
w_real[881] = 8'h51; w_imag[881] = 8'h62;
w_real[882] = 8'h52; w_imag[882] = 8'h61;
w_real[883] = 8'h53; w_imag[883] = 8'h61;
w_real[884] = 8'h53; w_imag[884] = 8'h60;
w_real[885] = 8'h54; w_imag[885] = 8'h60;
w_real[886] = 8'h54; w_imag[886] = 8'h5F;
w_real[887] = 8'h55; w_imag[887] = 8'h5F;
w_real[888] = 8'h55; w_imag[888] = 8'h5E;
w_real[889] = 8'h56; w_imag[889] = 8'h5E;
w_real[890] = 8'h57; w_imag[890] = 8'h5D;
w_real[891] = 8'h57; w_imag[891] = 8'h5D;
w_real[892] = 8'h58; w_imag[892] = 8'h5C;
w_real[893] = 8'h58; w_imag[893] = 8'h5C;
w_real[894] = 8'h59; w_imag[894] = 8'h5B;
w_real[895] = 8'h59; w_imag[895] = 8'h5B;
w_real[896] = 8'h5A; w_imag[896] = 8'h5A;
w_real[897] = 8'h5B; w_imag[897] = 8'h59;
w_real[898] = 8'h5B; w_imag[898] = 8'h59;
w_real[899] = 8'h5C; w_imag[899] = 8'h58;
w_real[900] = 8'h5C; w_imag[900] = 8'h58;
w_real[901] = 8'h5D; w_imag[901] = 8'h57;
w_real[902] = 8'h5D; w_imag[902] = 8'h57;
w_real[903] = 8'h5E; w_imag[903] = 8'h56;
w_real[904] = 8'h5E; w_imag[904] = 8'h55;
w_real[905] = 8'h5F; w_imag[905] = 8'h55;
w_real[906] = 8'h5F; w_imag[906] = 8'h54;
w_real[907] = 8'h60; w_imag[907] = 8'h54;
w_real[908] = 8'h60; w_imag[908] = 8'h53;
w_real[909] = 8'h61; w_imag[909] = 8'h53;
w_real[910] = 8'h61; w_imag[910] = 8'h52;
w_real[911] = 8'h62; w_imag[911] = 8'h51;
w_real[912] = 8'h62; w_imag[912] = 8'h51;
w_real[913] = 8'h63; w_imag[913] = 8'h50;
w_real[914] = 8'h63; w_imag[914] = 8'h4F;
w_real[915] = 8'h64; w_imag[915] = 8'h4F;
w_real[916] = 8'h64; w_imag[916] = 8'h4E;
w_real[917] = 8'h65; w_imag[917] = 8'h4E;
w_real[918] = 8'h65; w_imag[918] = 8'h4D;
w_real[919] = 8'h66; w_imag[919] = 8'h4C;
w_real[920] = 8'h66; w_imag[920] = 8'h4C;
w_real[921] = 8'h67; w_imag[921] = 8'h4B;
w_real[922] = 8'h67; w_imag[922] = 8'h4A;
w_real[923] = 8'h68; w_imag[923] = 8'h4A;
w_real[924] = 8'h68; w_imag[924] = 8'h49;
w_real[925] = 8'h69; w_imag[925] = 8'h49;
w_real[926] = 8'h69; w_imag[926] = 8'h48;
w_real[927] = 8'h69; w_imag[927] = 8'h47;
w_real[928] = 8'h6A; w_imag[928] = 8'h47;
w_real[929] = 8'h6A; w_imag[929] = 8'h46;
w_real[930] = 8'h6B; w_imag[930] = 8'h45;
w_real[931] = 8'h6B; w_imag[931] = 8'h45;
w_real[932] = 8'h6C; w_imag[932] = 8'h44;
w_real[933] = 8'h6C; w_imag[933] = 8'h43;
w_real[934] = 8'h6C; w_imag[934] = 8'h43;
w_real[935] = 8'h6D; w_imag[935] = 8'h42;
w_real[936] = 8'h6D; w_imag[936] = 8'h41;
w_real[937] = 8'h6E; w_imag[937] = 8'h41;
w_real[938] = 8'h6E; w_imag[938] = 8'h40;
w_real[939] = 8'h6E; w_imag[939] = 8'h3F;
w_real[940] = 8'h6F; w_imag[940] = 8'h3F;
w_real[941] = 8'h6F; w_imag[941] = 8'h3E;
w_real[942] = 8'h70; w_imag[942] = 8'h3D;
w_real[943] = 8'h70; w_imag[943] = 8'h3D;
w_real[944] = 8'h70; w_imag[944] = 8'h3C;
w_real[945] = 8'h71; w_imag[945] = 8'h3B;
w_real[946] = 8'h71; w_imag[946] = 8'h3A;
w_real[947] = 8'h71; w_imag[947] = 8'h3A;
w_real[948] = 8'h72; w_imag[948] = 8'h39;
w_real[949] = 8'h72; w_imag[949] = 8'h38;
w_real[950] = 8'h73; w_imag[950] = 8'h38;
w_real[951] = 8'h73; w_imag[951] = 8'h37;
w_real[952] = 8'h73; w_imag[952] = 8'h36;
w_real[953] = 8'h74; w_imag[953] = 8'h36;
w_real[954] = 8'h74; w_imag[954] = 8'h35;
w_real[955] = 8'h74; w_imag[955] = 8'h34;
w_real[956] = 8'h75; w_imag[956] = 8'h33;
w_real[957] = 8'h75; w_imag[957] = 8'h33;
w_real[958] = 8'h75; w_imag[958] = 8'h32;
w_real[959] = 8'h75; w_imag[959] = 8'h31;
w_real[960] = 8'h76; w_imag[960] = 8'h30;
w_real[961] = 8'h76; w_imag[961] = 8'h30;
w_real[962] = 8'h76; w_imag[962] = 8'h2F;
w_real[963] = 8'h77; w_imag[963] = 8'h2E;
w_real[964] = 8'h77; w_imag[964] = 8'h2E;
w_real[965] = 8'h77; w_imag[965] = 8'h2D;
w_real[966] = 8'h77; w_imag[966] = 8'h2C;
w_real[967] = 8'h78; w_imag[967] = 8'h2B;
w_real[968] = 8'h78; w_imag[968] = 8'h2B;
w_real[969] = 8'h78; w_imag[969] = 8'h2A;
w_real[970] = 8'h79; w_imag[970] = 8'h29;
w_real[971] = 8'h79; w_imag[971] = 8'h28;
w_real[972] = 8'h79; w_imag[972] = 8'h28;
w_real[973] = 8'h79; w_imag[973] = 8'h27;
w_real[974] = 8'h7A; w_imag[974] = 8'h26;
w_real[975] = 8'h7A; w_imag[975] = 8'h25;
w_real[976] = 8'h7A; w_imag[976] = 8'h25;
w_real[977] = 8'h7A; w_imag[977] = 8'h24;
w_real[978] = 8'h7A; w_imag[978] = 8'h23;
w_real[979] = 8'h7B; w_imag[979] = 8'h22;
w_real[980] = 8'h7B; w_imag[980] = 8'h22;
w_real[981] = 8'h7B; w_imag[981] = 8'h21;
w_real[982] = 8'h7B; w_imag[982] = 8'h20;
w_real[983] = 8'h7B; w_imag[983] = 8'h1F;
w_real[984] = 8'h7C; w_imag[984] = 8'h1F;
w_real[985] = 8'h7C; w_imag[985] = 8'h1E;
w_real[986] = 8'h7C; w_imag[986] = 8'h1D;
w_real[987] = 8'h7C; w_imag[987] = 8'h1C;
w_real[988] = 8'h7C; w_imag[988] = 8'h1C;
w_real[989] = 8'h7D; w_imag[989] = 8'h1B;
w_real[990] = 8'h7D; w_imag[990] = 8'h1A;
w_real[991] = 8'h7D; w_imag[991] = 8'h19;
w_real[992] = 8'h7D; w_imag[992] = 8'h18;
w_real[993] = 8'h7D; w_imag[993] = 8'h18;
w_real[994] = 8'h7D; w_imag[994] = 8'h17;
w_real[995] = 8'h7D; w_imag[995] = 8'h16;
w_real[996] = 8'h7E; w_imag[996] = 8'h15;
w_real[997] = 8'h7E; w_imag[997] = 8'h15;
w_real[998] = 8'h7E; w_imag[998] = 8'h14;
w_real[999] = 8'h7E; w_imag[999] = 8'h13;
w_real[1000] = 8'h7E; w_imag[1000] = 8'h12;
w_real[1001] = 8'h7E; w_imag[1001] = 8'h12;
w_real[1002] = 8'h7E; w_imag[1002] = 8'h11;
w_real[1003] = 8'h7E; w_imag[1003] = 8'h10;
w_real[1004] = 8'h7F; w_imag[1004] = 8'h0F;
w_real[1005] = 8'h7F; w_imag[1005] = 8'h0E;
w_real[1006] = 8'h7F; w_imag[1006] = 8'h0E;
w_real[1007] = 8'h7F; w_imag[1007] = 8'h0D;
w_real[1008] = 8'h7F; w_imag[1008] = 8'h0C;
w_real[1009] = 8'h7F; w_imag[1009] = 8'h0B;
w_real[1010] = 8'h7F; w_imag[1010] = 8'h0A;
w_real[1011] = 8'h7F; w_imag[1011] = 8'h0A;
w_real[1012] = 8'h7F; w_imag[1012] = 8'h09;
w_real[1013] = 8'h7F; w_imag[1013] = 8'h08;
w_real[1014] = 8'h7F; w_imag[1014] = 8'h07;
w_real[1015] = 8'h7F; w_imag[1015] = 8'h07;
w_real[1016] = 8'h7F; w_imag[1016] = 8'h06;
w_real[1017] = 8'h7F; w_imag[1017] = 8'h05;
w_real[1018] = 8'h7F; w_imag[1018] = 8'h04;
w_real[1019] = 8'h7F; w_imag[1019] = 8'h03;
w_real[1020] = 8'h7F; w_imag[1020] = 8'h03;
w_real[1021] = 8'h7F; w_imag[1021] = 8'h02;
w_real[1022] = 8'h7F; w_imag[1022] = 8'h01;
w_real[1023] = 8'h7F; w_imag[1023] = 8'h00;
