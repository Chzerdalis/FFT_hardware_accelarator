gen_input_real[0] = 24'sd0;
gen_input_real[4] = 24'sd2047;
gen_input_real[8] = -24'sd410;
gen_input_real[12] = -24'sd1505;
gen_input_real[1] = 24'sd560;
gen_input_real[5] = 24'sd1135;
gen_input_real[9] = -24'sd728;
gen_input_real[13] = -24'sd958;
gen_input_real[2] = 24'sd958;
gen_input_real[6] = 24'sd728;
gen_input_real[10] = -24'sd1135;
gen_input_real[14] = -24'sd560;
gen_input_real[3] = 24'sd1505;
gen_input_real[7] = 24'sd410;
gen_input_real[11] = -24'sd2047;
gen_input_real[15] = 24'sd0;
