0 0
0 -17
0 -28
0 -15
0 -5
0 -43
0 -50
1 -59
1 -54
1 -59
1 -57
2 -65
2 -68
3 -77
4 -107
5 -109
5 -103
5 -110
6 -109
8 -153
9 -151
9 -148
10 -156
11 -158
12 -172
12 -162
15 -191
15 -189
16 -190
18 -206
19 -207
21 -225
22 -228
26 -258
26 -256
26 -250
30 -270
31 -274
30 -261
35 -295
38 -308
51 -409
41 -316
59 -447
44 -328
45 -328
46 -329
48 -336
52 -356
54 -359
57 -373
60 -382
62 -388
67 -409
65 -393
72 -426
74 -427
81 -461
77 -433
87 -479
92 -499
208 -1103
208 -1084
84 -429
91 -458
99 -492
106 -518
107 -517
108 -513
117 -546
122 -561
128 -580
142 -636
408 -1792
113 -490
126 -538
138 -582
141 -586
148 -609
153 -619
163 -652
165 -652
166 -648
173 -667
180 -683
183 -686
187 -693
206 -754
203 -736
210 -751
213 -754
222 -776
230 -794
237 -811
245 -826
253 -844
261 -861
274 -896
280 -903
289 -922
305 -962
325 -1018
338 -1046
364 -1113
379 -1147
404 -1212
454 -1349
557 -1636
2346 -6821
228 -657
464 -1324
2517 -7104
55 -153
224 -622
300 -824
358 -974
410 -1103
488 -1300
653 -1725
3481 -9107
-46 119
180 -464
265 -675
314 -794
351 -879
383 -950
404 -994
429 -1045
448 -1082
470 -1124
501 -1189
515 -1213
533 -1245
559 -1294
585 -1343
619 -1409
650 -1466
681 -1523
719 -1596
772 -1699
838 -1831
948 -2055
1145 -2460
1611 -3434
8596 -18175
-616 1293
98 -205
324 -670
456 -934
536 -1090
613 -1237
664 -1331
716 -1423
779 -1537
833 -1630
884 -1718
951 -1834
1021 -1953
1112 -2111
1211 -2283
1344 -2516
1564 -2905
1933 -3564
2927 -5356
15812 -28729
-1925 3473
-344 616
152 -271
413 -729
572 -1003
706 -1229
799 -1380
893 -1532
979 -1669
1060 -1794
1141 -1918
1227 -2047
1319 -2185
1401 -2306
1522 -2487
1634 -2653
1763 -2843
1941 -3108
2156 -3429
2461 -3886
2935 -4604
3730 -5811
5854 -9059
30211 -46439
-4928 7524
-1268 1923
-121 183
492 -737
917 -1364
1262 -1864
1628 -2389
2002 -2918
2476 -3585
3179 -4573
4380 -6260
7421 -10537
40540 -57189
-8559 11996
-3122 4347
-1465 2027
-671 923
-160 218
193 -262
526 -709
752 -1008
971 -1293
1194 -1580
1400 -1840
1584 -2068
1820 -2362
2043 -2635
2290 -2934
2575 -3279
2941 -3722
3349 -4211
3907 -4882
4653 -5777
5840 -7206
7992 -9800
13535 -16493
68715 -83207
-17288 20804
-6534 7814
-3426 4071
-1915 2262
-982 1153
-283 330
210 -243
671 -773
1059 -1213
1421 -1617
1754 -1983
2103 -2364
2470 -2759
2847 -3160
3234 -3568
3655 -4008
4155 -4529
4736 -5130
5407 -5820
6193 -6625
7216 -7673
8517 -9001
10355 -10876
13112 -13687
17936 -18609
29335 -30249
122667 -125716
-23805 24247
8062 -8161
109875 -110551
-46973 46973
-22558 22420
-15253 15067
-11538 11327
-9214 8991
-7561 7332
-6325 6096
-5331 5107
-4488 4273
-3748 3546
-3077 2894
-2411 2253
-1746 1622
-1026 947
-197 181
792 -723
2093 -1897
4082 -3677
7589 -6794
16364 -14559
88755 -78481
-36742 32288
-17009 14855
-11609 10077
-9091 7842
-7561 6482
-6537 5569
-5763 4880
-5201 4376
-4717 3944
-4313 3584
-3977 3284
-3664 3007
-3389 2764
-3129 2536
-2867 2309
-2686 2150
-2463 1959
-2238 1769
-2037 1600
-1807 1410
-1582 1226
-1312 1011
-1042 798
-731 556
-375 283
64 -48
654 -488
1482 -1099
2690 -1982
4916 -3599
10391 -7559
51717 -37381
-25029 17974
-11330 8084
-7681 5445
-5991 4219
-4984 3487
-4302 2990
-3763 2599
-3353 2300
-3026 2062
-2714 1838
-2449 1647
-2202 1471
-1964 1304
-1734 1143
-1517 993
-1258 818
-966 624
-701 450
-363 231
-6 4
471 -296
1082 -676
1997 -1239
3524 -2172
7149 -4375
31457 -19118
-15621 9428
-6038 3619
-3261 1941
-1578 932
-123 72
1732 -1009
5249 -3038
25998 -14939
-13173 7516
-3744 2121
1278 -719
20800 -11615
-14861 8239
-6202 3413
-2769 1513
1171 -635
18809 -10127
-11295 6037
11166 -5924
-18225 9598
-10676 5581
-8446 4382
-7243 3729
-6429 3285
-5870 2977
-5416 2726
-5042 2518
-4732 2345
-4434 2181
-4148 2024
-3906 1891
-3615 1737
-3262 1555
-2817 1332
-2123 996
-583 271
8872 -4097
-11042 5057
-6533 2968
-5384 2426
-4816 2152
-4448 1971
-4193 1843
-4016 1751
-3845 1662
-3696 1584
-3561 1513
-3427 1444
-3283 1371
-3176 1315
-3046 1251
-2885 1174
-2670 1077
-2405 962
-2002 793
-1097 431
4007 -1559
-7052 2720
-4206 1607
-3246 1229
-2238 839
2153 -800
-7245 2667
-4838 1764
-4197 1516
-3859 1380
-3653 1294
-3467 1216
-3336 1159
-3194 1098
-3017 1027
-2755 929
-2258 753
492 -162
-5689 1860
-4123 1334
-3698 1184
-3509 1111
-3361 1053
-3271 1014
-3169 972
-3072 931
-2960 888
-2810 833
-2491 730
-842 244
-4688 1344
-3665 1038
-3438 962
-3264 903
-3195 873
-3149 850
-3096 826
-3064 807
-3036 790
-2999 770
-2970 753
-2945 737
-2931 724
-2899 707
-2901 698
-2875 682
-2847 666
-2854 659
-2854 650
-2815 632
-2793 618
-2787 608
-2769 595
-2773 587
-2731 569
-2749 564
-2723 550
-2725 542
-2713 531
-2708 521
-2691 509
-2679 498
-2687 491
-2661 478
-2656 469
-2646 459
-2662 453
-2639 441
-2625 430
-2639 424
-2621 413
-2614 404
-2603 394
-2598 385
-2608 378
-2577 366
-2580 358
-2582 350
-2577 342
-2559 331
-2578 326
-2564 316
-2556 307
-2570 301
-2548 290
-2549 282
-2534 273
-2516 263
-2534 257
-2516 247
-2524 240
-2502 230
-2494 222
-2517 216
-2509 208
-2506 200
-2488 191
-2511 185
-2508 177
-2499 168
-2513 162
-2484 152
-2497 145
-2495 137
-2505 130
-2506 123
-2479 114
-2479 106
-2489 99
-2478 91
-2479 83
-2465 75
-2460 67
-2478 60
-2471 53
-2462 45
-2501 38
-2492 30
-2470 22
-2474 15
-2485 7
-2486 0
-2485 -7
-2474 -15
-2470 -22
-2492 -30
-2501 -38
-2462 -45
-2471 -53
-2478 -60
-2460 -67
-2465 -75
-2479 -83
-2478 -91
-2489 -99
-2479 -106
-2479 -114
-2506 -123
-2505 -130
-2495 -137
-2497 -145
-2484 -152
-2513 -162
-2499 -168
-2508 -177
-2511 -185
-2488 -191
-2506 -200
-2509 -208
-2517 -216
-2494 -222
-2502 -230
-2524 -240
-2516 -247
-2534 -257
-2516 -263
-2534 -273
-2549 -282
-2548 -290
-2570 -301
-2556 -307
-2564 -316
-2578 -326
-2559 -331
-2577 -342
-2582 -350
-2580 -358
-2577 -366
-2608 -378
-2598 -385
-2603 -394
-2614 -404
-2621 -413
-2639 -424
-2625 -430
-2639 -441
-2662 -453
-2646 -459
-2656 -469
-2661 -478
-2687 -491
-2679 -498
-2691 -509
-2708 -521
-2713 -531
-2725 -542
-2723 -550
-2749 -564
-2731 -569
-2773 -587
-2769 -595
-2787 -608
-2793 -618
-2815 -632
-2854 -650
-2854 -659
-2847 -666
-2875 -682
-2901 -698
-2899 -707
-2931 -724
-2945 -737
-2970 -753
-2999 -770
-3036 -790
-3064 -807
-3096 -826
-3149 -850
-3195 -873
-3264 -903
-3438 -962
-3665 -1038
-4688 -1344
-842 -244
-2491 -730
-2810 -833
-2960 -888
-3072 -931
-3169 -972
-3271 -1014
-3361 -1053
-3509 -1111
-3698 -1184
-4123 -1334
-5689 -1860
492 162
-2258 -753
-2755 -929
-3017 -1027
-3194 -1098
-3336 -1159
-3467 -1216
-3653 -1294
-3859 -1380
-4197 -1516
-4838 -1764
-7245 -2667
2153 800
-2238 -839
-3246 -1229
-4206 -1607
-7052 -2720
4007 1559
-1097 -431
-2002 -793
-2405 -962
-2670 -1077
-2885 -1174
-3046 -1251
-3176 -1315
-3283 -1371
-3427 -1444
-3561 -1513
-3696 -1584
-3845 -1662
-4016 -1751
-4193 -1843
-4448 -1971
-4816 -2152
-5384 -2426
-6533 -2968
-11042 -5057
8872 4097
-583 -271
-2123 -996
-2817 -1332
-3262 -1555
-3615 -1737
-3906 -1891
-4148 -2024
-4434 -2181
-4732 -2345
-5042 -2518
-5416 -2726
-5870 -2977
-6429 -3285
-7243 -3729
-8446 -4382
-10676 -5581
-18225 -9598
11166 5924
-11295 -6037
18809 10127
1171 635
-2769 -1513
-6202 -3413
-14861 -8239
20800 11615
1278 719
-3744 -2121
-13173 -7516
25998 14939
5249 3038
1732 1009
-123 -72
-1578 -932
-3261 -1941
-6038 -3619
-15621 -9428
31457 19118
7149 4375
3524 2172
1997 1239
1082 676
471 296
-6 -4
-363 -231
-701 -450
-966 -624
-1258 -818
-1517 -993
-1734 -1143
-1964 -1304
-2202 -1471
-2449 -1647
-2714 -1838
-3026 -2062
-3353 -2300
-3763 -2599
-4302 -2990
-4984 -3487
-5991 -4219
-7681 -5445
-11330 -8084
-25029 -17974
51717 37381
10391 7559
4916 3599
2690 1982
1482 1099
654 488
64 48
-375 -283
-731 -556
-1042 -798
-1312 -1011
-1582 -1226
-1807 -1410
-2037 -1600
-2238 -1769
-2463 -1959
-2686 -2150
-2867 -2309
-3129 -2536
-3389 -2764
-3664 -3007
-3977 -3284
-4313 -3584
-4717 -3944
-5201 -4376
-5763 -4880
-6537 -5569
-7561 -6482
-9091 -7842
-11609 -10077
-17009 -14855
-36742 -32288
88755 78481
16364 14559
7589 6794
4082 3677
2093 1897
792 723
-197 -181
-1026 -947
-1746 -1622
-2411 -2253
-3077 -2894
-3748 -3546
-4488 -4273
-5331 -5107
-6325 -6096
-7561 -7332
-9214 -8991
-11538 -11327
-15253 -15067
-22558 -22420
-46973 -46973
109875 110551
8062 8161
-23805 -24247
122667 125716
29335 30249
17936 18609
13112 13687
10355 10876
8517 9001
7216 7673
6193 6625
5407 5820
4736 5130
4155 4529
3655 4008
3234 3568
2847 3160
2470 2759
2103 2364
1754 1983
1421 1617
1059 1213
671 773
210 243
-283 -330
-982 -1153
-1915 -2262
-3426 -4071
-6534 -7814
-17288 -20804
68715 83207
13535 16493
7992 9800
5840 7206
4653 5777
3907 4882
3349 4211
2941 3722
2575 3279
2290 2934
2043 2635
1820 2362
1584 2068
1400 1840
1194 1580
971 1293
752 1008
526 709
193 262
-160 -218
-671 -923
-1465 -2027
-3122 -4347
-8559 -11996
40540 57189
7421 10537
4380 6260
3179 4573
2476 3585
2002 2918
1628 2389
1262 1864
917 1364
492 737
-121 -183
-1268 -1923
-4928 -7524
30211 46439
5854 9059
3730 5811
2935 4604
2461 3886
2156 3429
1941 3108
1763 2843
1634 2653
1522 2487
1401 2306
1319 2185
1227 2047
1141 1918
1060 1794
979 1669
893 1532
799 1380
706 1229
572 1003
413 729
152 271
-344 -616
-1925 -3473
15812 28729
2927 5356
1933 3564
1564 2905
1344 2516
1211 2283
1112 2111
1021 1953
951 1834
884 1718
833 1630
779 1537
716 1423
664 1331
613 1237
536 1090
456 934
324 670
98 205
-616 -1293
8596 18175
1611 3434
1145 2460
948 2055
838 1831
772 1699
719 1596
681 1523
650 1466
619 1409
585 1343
559 1294
533 1245
515 1213
501 1189
470 1124
448 1082
429 1045
404 994
383 950
351 879
314 794
265 675
180 464
-46 -119
3481 9107
653 1725
488 1300
410 1103
358 974
300 824
224 622
55 153
2517 7104
464 1324
228 657
2346 6821
557 1636
454 1349
404 1212
379 1147
364 1113
338 1046
325 1018
305 962
289 922
280 903
274 896
261 861
253 844
245 826
237 811
230 794
222 776
213 754
210 751
203 736
206 754
187 693
183 686
180 683
173 667
166 648
165 652
163 652
153 619
148 609
141 586
138 582
126 538
113 490
408 1792
142 636
128 580
122 561
117 546
108 513
107 517
106 518
99 492
91 458
84 429
208 1084
208 1103
92 499
87 479
77 433
81 461
74 427
72 426
65 393
67 409
62 388
60 382
57 373
54 359
52 356
48 336
46 329
45 328
44 328
59 447
41 316
51 409
38 308
35 295
30 261
31 274
30 270
26 250
26 256
26 258
22 228
21 225
19 207
18 206
16 190
15 189
15 191
12 162
12 172
11 158
10 156
9 148
9 151
8 153
6 109
5 110
5 103
5 109
4 107
3 77
2 68
2 65
1 57
1 59
1 54
1 59
0 50
0 43
0 5
0 15
0 28
0 17
