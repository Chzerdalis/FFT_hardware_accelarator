0 0
0 0
0 -7
0 0
0 14
0 -5
0 0
0 3
0 -2
0 -4
0 10
0 -26
0 11
0 -8
0 -10
0 3
0 -9
1 -21
1 -19
1 -31
2 -37
1 -25
1 -17
0 -1
1 -24
1 -21
1 -22
2 -31
3 -36
2 -25
3 -42
2 -22
1 -13
3 -31
4 -40
1 -15
1 -16
3 -33
3 -29
4 -35
4 -34
7 -56
6 -52
7 -54
6 -46
5 -37
5 -40
6 -43
7 -47
3 -20
7 -48
5 -37
8 -54
10 -61
9 -57
9 -53
10 -58
11 -62
7 -42
10 -59
10 -54
27 -144
25 -134
9 -48
8 -42
11 -56
10 -51
14 -70
12 -60
13 -63
15 -71
15 -71
18 -84
51 -224
17 -74
13 -58
13 -58
15 -63
18 -77
21 -88
19 -77
23 -94
24 -95
23 -89
20 -78
18 -69
20 -74
29 -109
23 -83
29 -104
28 -100
28 -100
30 -105
25 -85
29 -100
26 -89
36 -121
31 -103
34 -109
35 -112
34 -109
36 -113
41 -128
54 -165
51 -155
54 -163
59 -177
66 -196
288 -839
35 -101
56 -161
315 -890
5 -14
26 -73
37 -103
44 -119
52 -141
62 -165
82 -217
432 -1131
0 0
25 -66
32 -81
37 -95
48 -121
56 -140
49 -121
48 -117
55 -135
55 -133
64 -152
61 -143
70 -164
59 -137
65 -150
80 -183
79 -179
86 -192
84 -186
96 -212
101 -221
115 -249
141 -303
210 -449
1068 -2258
-69 144
15 -33
37 -76
65 -134
63 -129
78 -157
77 -154
87 -173
101 -200
115 -226
109 -213
121 -234
127 -244
141 -268
166 -313
173 -324
200 -372
242 -447
371 -680
1971 -3581
-229 414
-43 77
36 -64
61 -108
71 -125
79 -138
102 -177
117 -200
120 -204
130 -220
132 -222
157 -263
165 -274
170 -281
191 -313
200 -326
212 -342
255 -409
266 -424
314 -496
359 -563
449 -700
729 -1128
3728 -5730
-616 941
-168 255
-15 22
55 -82
124 -184
156 -231
192 -283
241 -351
306 -443
380 -547
558 -798
926 -1314
5027 -7092
-1053 1477
-389 542
-156 217
-76 104
-26 36
9 -12
75 -102
94 -126
119 -159
156 -207
185 -243
193 -252
224 -290
250 -322
274 -351
320 -407
378 -479
423 -532
497 -621
580 -720
733 -905
995 -1220
1674 -2040
8514 -10310
-2147 2584
-794 949
-397 472
-240 283
-131 154
-19 22
9 -11
83 -95
128 -147
180 -205
205 -232
256 -288
310 -346
362 -402
401 -442
453 -496
506 -551
590 -639
675 -727
777 -832
909 -967
1065 -1125
1275 -1339
1635 -1707
2220 -2303
3626 -3739
15185 -15562
-2950 3005
988 -1000
13609 -13693
-5822 5822
-2785 2768
-1886 1863
-1422 1396
-1138 1110
-933 904
-789 760
-661 633
-550 523
-480 454
-389 366
-291 272
-225 209
-133 123
-15 14
105 -96
254 -230
532 -479
953 -853
2027 -1803
11007 -9733
-4539 3989
-2108 1841
-1412 1226
-1156 997
-953 817
-814 693
-704 596
-657 553
-587 491
-548 455
-477 393
-457 375
-422 344
-369 299
-338 272
-335 268
-312 248
-269 213
-262 205
-225 176
-190 147
-161 124
-127 97
-85 64
-49 37
6 -4
89 -66
204 -151
348 -256
631 -462
1289 -937
6401 -4627
-3102 2227
-1409 1005
-923 654
-751 528
-621 434
-540 375
-464 321
-419 287
-365 249
-330 223
-288 193
-259 173
-238 158
-221 145
-218 142
-175 114
-104 67
-101 64
-26 16
-25 15
76 -48
118 -74
229 -142
430 -265
862 -527
3897 -2368
-1951 1177
-755 452
-421 250
-187 110
-26 15
221 -129
656 -380
3217 -1848
-1615 922
-466 264
156 -88
2574 -1437
-1854 1027
-779 428
-347 189
149 -81
2336 -1257
-1390 743
1377 -731
-2245 1182
-1332 696
-1053 546
-913 470
-778 397
-732 371
-675 340
-647 323
-590 292
-552 271
-513 250
-492 238
-452 217
-406 193
-356 168
-249 117
-79 36
1098 -507
-1357 621
-825 374
-670 302
-610 272
-533 236
-500 220
-505 220
-484 209
-473 202
-444 189
-409 172
-408 170
-407 168
-388 159
-359 146
-320 129
-313 125
-246 97
-137 54
501 -195
-885 341
-512 196
-403 152
-259 97
245 -91
-884 325
-606 221
-525 189
-477 170
-458 162
-438 153
-403 140
-398 137
-379 129
-334 112
-284 95
67 -22
-689 225
-505 163
-469 150
-447 141
-412 129
-397 123
-374 114
-387 117
-355 106
-355 105
-305 89
-108 31
-581 166
-445 126
-427 119
-405 112
-409 112
-375 101
-395 105
-370 97
-385 100
-361 92
-359 91
-355 88
-361 89
-366 89
-376 90
-344 81
-359 84
-369 85
-358 81
-361 81
-342 75
-338 73
-358 76
-331 70
-336 70
-344 70
-337 68
-348 69
-317 62
-342 65
-323 61
-331 61
-328 60
-324 58
-348 61
-332 57
-335 57
-333 55
-329 53
-329 53
-326 51
-314 48
-321 48
-320 47
-332 48
-320 45
-317 44
-323 43
-310 41
-327 42
-338 42
-322 39
-323 38
-305 35
-310 35
-309 34
-329 35
-307 32
-334 34
-298 29
-323 30
-319 29
-298 26
-308 26
-313 25
-297 23
-306 23
-330 24
-300 21
-309 20
-334 21
-299 18
-316 18
-285 15
-308 16
-312 15
-316 14
-309 13
-312 12
-317 11
-314 10
-308 9
-312 8
-310 7
-303 6
-310 5
-320 4
-340 4
-313 2
-321 1
-305 0
-308 0
-305 0
-321 -1
-313 -2
-340 -4
-320 -4
-310 -5
-303 -6
-310 -7
-312 -8
-308 -9
-314 -10
-317 -11
-312 -12
-309 -13
-316 -14
-312 -15
-308 -16
-285 -15
-316 -18
-299 -18
-334 -21
-309 -20
-300 -21
-330 -24
-306 -23
-297 -23
-313 -25
-308 -26
-298 -26
-319 -29
-323 -30
-298 -29
-334 -34
-307 -32
-329 -35
-309 -34
-310 -35
-305 -35
-323 -38
-322 -39
-338 -42
-327 -42
-310 -41
-323 -43
-317 -44
-320 -45
-332 -48
-320 -47
-321 -48
-314 -48
-326 -51
-329 -53
-329 -53
-333 -55
-335 -57
-332 -57
-348 -61
-324 -58
-328 -60
-331 -61
-323 -61
-342 -65
-317 -62
-348 -69
-337 -68
-344 -70
-336 -70
-331 -70
-358 -76
-338 -73
-342 -75
-361 -81
-358 -81
-369 -85
-359 -84
-344 -81
-376 -90
-366 -89
-361 -89
-355 -88
-359 -91
-361 -92
-385 -100
-370 -97
-395 -105
-375 -101
-409 -112
-405 -112
-427 -119
-445 -126
-581 -166
-108 -31
-305 -89
-355 -105
-355 -106
-387 -117
-374 -114
-397 -123
-412 -129
-447 -141
-469 -150
-505 -163
-689 -225
67 22
-284 -95
-334 -112
-379 -129
-398 -137
-403 -140
-438 -153
-458 -162
-477 -170
-525 -189
-606 -221
-884 -325
245 91
-259 -97
-403 -152
-512 -196
-885 -341
501 195
-137 -54
-246 -97
-313 -125
-320 -129
-359 -146
-388 -159
-407 -168
-408 -170
-409 -172
-444 -189
-473 -202
-484 -209
-505 -220
-500 -220
-533 -236
-610 -272
-670 -302
-825 -374
-1357 -621
1098 507
-79 -36
-249 -117
-356 -168
-406 -193
-452 -217
-492 -238
-513 -250
-552 -271
-590 -292
-647 -323
-675 -340
-732 -371
-778 -397
-913 -470
-1053 -546
-1332 -696
-2245 -1182
1377 731
-1390 -743
2336 1257
149 81
-347 -189
-779 -428
-1854 -1027
2574 1437
156 88
-466 -264
-1615 -922
3217 1848
656 380
221 129
-26 -15
-187 -110
-421 -250
-755 -452
-1951 -1177
3897 2368
862 527
430 265
229 142
118 74
76 48
-25 -15
-26 -16
-101 -64
-104 -67
-175 -114
-218 -142
-221 -145
-238 -158
-259 -173
-288 -193
-330 -223
-365 -249
-419 -287
-464 -321
-540 -375
-621 -434
-751 -528
-923 -654
-1409 -1005
-3102 -2227
6401 4627
1289 937
631 462
348 256
204 151
89 66
6 4
-49 -37
-85 -64
-127 -97
-161 -124
-190 -147
-225 -176
-262 -205
-269 -213
-312 -248
-335 -268
-338 -272
-369 -299
-422 -344
-457 -375
-477 -393
-548 -455
-587 -491
-657 -553
-704 -596
-814 -693
-953 -817
-1156 -997
-1412 -1226
-2108 -1841
-4539 -3989
11007 9733
2027 1803
953 853
532 479
254 230
105 96
-15 -14
-133 -123
-225 -209
-291 -272
-389 -366
-480 -454
-550 -523
-661 -633
-789 -760
-933 -904
-1138 -1110
-1422 -1396
-1886 -1863
-2785 -2768
-5822 -5822
13609 13693
988 1000
-2950 -3005
15185 15562
3626 3739
2220 2303
1635 1707
1275 1339
1065 1125
909 967
777 832
675 727
590 639
506 551
453 496
401 442
362 402
310 346
256 288
205 232
180 205
128 147
83 95
9 11
-19 -22
-131 -154
-240 -283
-397 -472
-794 -949
-2147 -2584
8514 10310
1674 2040
995 1220
733 905
580 720
497 621
423 532
378 479
320 407
274 351
250 322
224 290
193 252
185 243
156 207
119 159
94 126
75 102
9 12
-26 -36
-76 -104
-156 -217
-389 -542
-1053 -1477
5027 7092
926 1314
558 798
380 547
306 443
241 351
192 283
156 231
124 184
55 82
-15 -22
-168 -255
-616 -941
3728 5730
729 1128
449 700
359 563
314 496
266 424
255 409
212 342
200 326
191 313
170 281
165 274
157 263
132 222
130 220
120 204
117 200
102 177
79 138
71 125
61 108
36 64
-43 -77
-229 -414
1971 3581
371 680
242 447
200 372
173 324
166 313
141 268
127 244
121 234
109 213
115 226
101 200
87 173
77 154
78 157
63 129
65 134
37 76
15 33
-69 -144
1068 2258
210 449
141 303
115 249
101 221
96 212
84 186
86 192
79 179
80 183
65 150
59 137
70 164
61 143
64 152
55 133
55 135
48 117
49 121
56 140
48 121
37 95
32 81
25 66
0 0
432 1131
82 217
62 165
52 141
44 119
37 103
26 73
5 14
315 890
56 161
35 101
288 839
66 196
59 177
54 163
51 155
54 165
41 128
36 113
34 109
35 112
34 109
31 103
36 121
26 89
29 100
25 85
30 105
28 100
28 100
29 104
23 83
29 109
20 74
18 69
20 78
23 89
24 95
23 94
19 77
21 88
18 77
15 63
13 58
13 58
17 74
51 224
18 84
15 71
15 71
13 63
12 60
14 70
10 51
11 56
8 42
9 48
25 134
27 144
10 54
10 59
7 42
11 62
10 58
9 53
9 57
10 61
8 54
5 37
7 48
3 20
7 47
6 43
5 40
5 37
6 46
7 54
6 52
7 56
4 34
4 35
3 29
3 33
1 16
1 15
4 40
3 31
1 13
2 22
3 42
2 25
3 36
2 31
1 22
1 21
1 24
0 1
1 17
1 25
2 37
1 31
1 19
1 21
0 9
0 -3
0 10
0 8
0 -11
0 26
0 -10
0 4
0 2
0 -3
0 0
0 5
0 -14
0 0
0 7
0 0
