0 0
89 -1829
372 -3779
850 -5732
1906 -9586
2567 -10249
5558 -18325
5435 -15189
8187 -19765
12290 -25986
19761 -36971
59432 -99156
90962 -136135
13233 -17843
127164 -154950
67594 -74578
86234 -86234
103175 -93513
-41186 33800
-84880 62951
-55171 36864
-41104 24637
-19102 10210
-23477 11104
-40719 16866
-52311 18717
-42886 13009
-38632 9676
-38194 7597
-37046 5495
-36434 3588
-35839 1760
-35660 0
-35839 -1760
-36434 -3588
-37046 -5495
-38194 -7597
-38632 -9676
-42886 -13009
-52311 -18717
-40719 -16866
-23477 -11104
-19102 -10210
-41104 -24637
-55171 -36864
-84880 -62951
-41186 -33800
103175 93513
86234 86234
67594 74578
127164 154950
13233 17843
90962 136135
59432 99156
19761 36971
12290 25986
8187 19765
5435 15189
5558 18325
2567 10249
1906 9586
850 5732
372 3779
89 1829
