gen_input_real[0] = 24'sd0;
gen_input_real[64] = 24'sd2047;
gen_input_real[128] = -24'sd39;
gen_input_real[192] = -24'sd1326;
gen_input_real[16] = -24'sd4;
gen_input_real[80] = 24'sd735;
gen_input_real[144] = 24'sd41;
gen_input_real[208] = -24'sd552;
gen_input_real[32] = -24'sd68;
gen_input_real[96] = 24'sd471;
gen_input_real[160] = 24'sd261;
gen_input_real[224] = -24'sd287;
gen_input_real[48] = -24'sd616;
gen_input_real[112] = 24'sd67;
gen_input_real[176] = 24'sd875;
gen_input_real[240] = -24'sd3;
gen_input_real[4] = -24'sd942;
gen_input_real[68] = 24'sd123;
gen_input_real[132] = 24'sd1011;
gen_input_real[196] = -24'sd304;
gen_input_real[20] = -24'sd1142;
gen_input_real[84] = 24'sd459;
gen_input_real[148] = 24'sd1154;
gen_input_real[212] = -24'sd503;
gen_input_real[36] = -24'sd1065;
gen_input_real[100] = 24'sd348;
gen_input_real[164] = 24'sd1072;
gen_input_real[228] = -24'sd56;
gen_input_real[52] = -24'sd1103;
gen_input_real[116] = -24'sd191;
gen_input_real[180] = 24'sd872;
gen_input_real[244] = 24'sd321;
gen_input_real[8] = -24'sd382;
gen_input_real[72] = -24'sd397;
gen_input_real[136] = 24'sd4;
gen_input_real[200] = 24'sd461;
gen_input_real[24] = 24'sd53;
gen_input_real[88] = -24'sd561;
gen_input_real[152] = -24'sd15;
gen_input_real[216] = 24'sd831;
gen_input_real[40] = 24'sd51;
gen_input_real[104] = -24'sd1160;
gen_input_real[168] = 24'sd27;
gen_input_real[232] = 24'sd1140;
gen_input_real[56] = -24'sd329;
gen_input_real[120] = -24'sd755;
gen_input_real[184] = 24'sd634;
gen_input_real[248] = 24'sd486;
gen_input_real[12] = -24'sd725;
gen_input_real[76] = -24'sd492;
gen_input_real[140] = 24'sd576;
gen_input_real[204] = 24'sd449;
gen_input_real[28] = -24'sd279;
gen_input_real[92] = -24'sd212;
gen_input_real[156] = -24'sd66;
gen_input_real[220] = -24'sd30;
gen_input_real[44] = 24'sd423;
gen_input_real[108] = 24'sd104;
gen_input_real[172] = -24'sd786;
gen_input_real[236] = 24'sd54;
gen_input_real[60] = 24'sd1070;
gen_input_real[124] = -24'sd283;
gen_input_real[188] = -24'sd1035;
gen_input_real[252] = 24'sd338;
gen_input_real[1] = 24'sd604;
gen_input_real[65] = -24'sd307;
gen_input_real[129] = -24'sd135;
gen_input_real[193] = 24'sd305;
gen_input_real[17] = -24'sd15;
gen_input_real[81] = -24'sd288;
gen_input_real[145] = -24'sd44;
gen_input_real[209] = 24'sd302;
gen_input_real[33] = -24'sd19;
gen_input_real[97] = -24'sd285;
gen_input_real[161] = 24'sd234;
gen_input_real[225] = 24'sd157;
gen_input_real[49] = -24'sd325;
gen_input_real[113] = -24'sd40;
gen_input_real[177] = 24'sd155;
gen_input_real[241] = -24'sd58;
gen_input_real[5] = 24'sd85;
gen_input_real[69] = 24'sd239;
gen_input_real[133] = -24'sd181;
gen_input_real[197] = -24'sd425;
gen_input_real[21] = 24'sd183;
gen_input_real[85] = 24'sd470;
gen_input_real[149] = -24'sd219;
gen_input_real[213] = -24'sd403;
gen_input_real[37] = 24'sd253;
gen_input_real[101] = 24'sd332;
gen_input_real[165] = -24'sd269;
gen_input_real[229] = -24'sd106;
gen_input_real[53] = 24'sd311;
gen_input_real[117] = -24'sd417;
gen_input_real[181] = -24'sd288;
gen_input_real[245] = 24'sd888;
gen_input_real[9] = 24'sd185;
gen_input_real[73] = -24'sd920;
gen_input_real[137] = -24'sd86;
gen_input_real[201] = 24'sd665;
gen_input_real[25] = -24'sd120;
gen_input_real[89] = -24'sd422;
gen_input_real[153] = 24'sd418;
gen_input_real[217] = 24'sd206;
gen_input_real[41] = -24'sd442;
gen_input_real[105] = 24'sd75;
gen_input_real[169] = 24'sd38;
gen_input_real[233] = -24'sd417;
gen_input_real[57] = 24'sd390;
gen_input_real[121] = 24'sd640;
gen_input_real[185] = -24'sd408;
gen_input_real[249] = -24'sd592;
gen_input_real[13] = 24'sd186;
gen_input_real[77] = 24'sd367;
gen_input_real[141] = -24'sd257;
gen_input_real[205] = -24'sd50;
gen_input_real[29] = 24'sd647;
gen_input_real[93] = -24'sd314;
gen_input_real[157] = -24'sd844;
gen_input_real[221] = 24'sd500;
gen_input_real[45] = 24'sd649;
gen_input_real[109] = -24'sd350;
gen_input_real[173] = -24'sd359;
gen_input_real[237] = 24'sd111;
gen_input_real[61] = 24'sd252;
gen_input_real[125] = -24'sd2;
gen_input_real[189] = -24'sd227;
gen_input_real[253] = -24'sd107;
gen_input_real[2] = 24'sd107;
gen_input_real[66] = 24'sd227;
gen_input_real[130] = 24'sd2;
gen_input_real[194] = -24'sd252;
gen_input_real[18] = -24'sd111;
gen_input_real[82] = 24'sd359;
gen_input_real[146] = 24'sd350;
gen_input_real[210] = -24'sd649;
gen_input_real[34] = -24'sd500;
gen_input_real[98] = 24'sd844;
gen_input_real[162] = 24'sd314;
gen_input_real[226] = -24'sd647;
gen_input_real[50] = 24'sd50;
gen_input_real[114] = 24'sd257;
gen_input_real[178] = -24'sd367;
gen_input_real[242] = -24'sd186;
gen_input_real[6] = 24'sd592;
gen_input_real[70] = 24'sd408;
gen_input_real[134] = -24'sd640;
gen_input_real[198] = -24'sd390;
gen_input_real[22] = 24'sd417;
gen_input_real[86] = -24'sd38;
gen_input_real[150] = -24'sd75;
gen_input_real[214] = 24'sd442;
gen_input_real[38] = -24'sd206;
gen_input_real[102] = -24'sd418;
gen_input_real[166] = 24'sd422;
gen_input_real[230] = 24'sd120;
gen_input_real[54] = -24'sd665;
gen_input_real[118] = 24'sd86;
gen_input_real[182] = 24'sd920;
gen_input_real[246] = -24'sd185;
gen_input_real[10] = -24'sd888;
gen_input_real[74] = 24'sd288;
gen_input_real[138] = 24'sd417;
gen_input_real[202] = -24'sd311;
gen_input_real[26] = 24'sd106;
gen_input_real[90] = 24'sd269;
gen_input_real[154] = -24'sd332;
gen_input_real[218] = -24'sd253;
gen_input_real[42] = 24'sd403;
gen_input_real[106] = 24'sd219;
gen_input_real[170] = -24'sd470;
gen_input_real[234] = -24'sd183;
gen_input_real[58] = 24'sd425;
gen_input_real[122] = 24'sd181;
gen_input_real[186] = -24'sd239;
gen_input_real[250] = -24'sd85;
gen_input_real[14] = 24'sd58;
gen_input_real[78] = -24'sd155;
gen_input_real[142] = 24'sd40;
gen_input_real[206] = 24'sd325;
gen_input_real[30] = -24'sd157;
gen_input_real[94] = -24'sd234;
gen_input_real[158] = 24'sd285;
gen_input_real[222] = 24'sd19;
gen_input_real[46] = -24'sd302;
gen_input_real[110] = 24'sd44;
gen_input_real[174] = 24'sd288;
gen_input_real[238] = 24'sd15;
gen_input_real[62] = -24'sd305;
gen_input_real[126] = 24'sd135;
gen_input_real[190] = 24'sd307;
gen_input_real[254] = -24'sd604;
gen_input_real[3] = -24'sd338;
gen_input_real[67] = 24'sd1035;
gen_input_real[131] = 24'sd283;
gen_input_real[195] = -24'sd1070;
gen_input_real[19] = -24'sd54;
gen_input_real[83] = 24'sd786;
gen_input_real[147] = -24'sd104;
gen_input_real[211] = -24'sd423;
gen_input_real[35] = 24'sd30;
gen_input_real[99] = 24'sd66;
gen_input_real[163] = 24'sd212;
gen_input_real[227] = 24'sd279;
gen_input_real[51] = -24'sd449;
gen_input_real[115] = -24'sd576;
gen_input_real[179] = 24'sd492;
gen_input_real[243] = 24'sd725;
gen_input_real[7] = -24'sd486;
gen_input_real[71] = -24'sd634;
gen_input_real[135] = 24'sd755;
gen_input_real[199] = 24'sd329;
gen_input_real[23] = -24'sd1140;
gen_input_real[87] = -24'sd27;
gen_input_real[151] = 24'sd1160;
gen_input_real[215] = -24'sd51;
gen_input_real[39] = -24'sd831;
gen_input_real[103] = 24'sd15;
gen_input_real[167] = 24'sd561;
gen_input_real[231] = -24'sd53;
gen_input_real[55] = -24'sd461;
gen_input_real[119] = -24'sd4;
gen_input_real[183] = 24'sd397;
gen_input_real[247] = 24'sd382;
gen_input_real[11] = -24'sd321;
gen_input_real[75] = -24'sd872;
gen_input_real[139] = 24'sd191;
gen_input_real[203] = 24'sd1103;
gen_input_real[27] = 24'sd56;
gen_input_real[91] = -24'sd1072;
gen_input_real[155] = -24'sd348;
gen_input_real[219] = 24'sd1065;
gen_input_real[43] = 24'sd503;
gen_input_real[107] = -24'sd1154;
gen_input_real[171] = -24'sd459;
gen_input_real[235] = 24'sd1142;
gen_input_real[59] = 24'sd304;
gen_input_real[123] = -24'sd1011;
gen_input_real[187] = -24'sd123;
gen_input_real[251] = 24'sd942;
gen_input_real[15] = 24'sd3;
gen_input_real[79] = -24'sd875;
gen_input_real[143] = -24'sd67;
gen_input_real[207] = 24'sd616;
gen_input_real[31] = 24'sd287;
gen_input_real[95] = -24'sd261;
gen_input_real[159] = -24'sd471;
gen_input_real[223] = 24'sd68;
gen_input_real[47] = 24'sd552;
gen_input_real[111] = -24'sd41;
gen_input_real[175] = -24'sd735;
gen_input_real[239] = 24'sd4;
gen_input_real[63] = 24'sd1326;
gen_input_real[127] = 24'sd39;
gen_input_real[191] = -24'sd2047;
gen_input_real[255] = 24'sd0;
