0 0
0 -10
0 -14
0 -6
1 -21
1 -26
1 -25
1 -16
3 -32
4 -44
3 -30
5 -42
8 -59
6 -39
9 -56
11 -59
17 -90
13 -65
14 -64
20 -87
35 -142
22 -86
23 -84
30 -103
66 -218
28 -91
36 -110
39 -115
47 -132
51 -139
58 -151
64 -162
68 -164
86 -201
105 -238
145 -317
606 -1282
11 -23
75 -150
112 -216
166 -311
615 -1118
91 -160
680 -1168
-31 51
60 -98
98 -155
142 -219
173 -260
227 -331
285 -405
428 -593
1711 -2307
-146 191
116 -148
236 -295
345 -420
478 -569
683 -792
1117 -1263
3925 -4331
2943 -3168
2039 -2141
-1765 1809
-906 906
-597 582
-411 391
-287 266
-168 153
-56 50
76 -66
304 -255
791 -649
4419 -3536
-2022 1578
-902 686
-536 397
-226 163
1116 -786
-1166 800
-695 464
-538 350
-450 285
-382 235
-291 174
-170 99
476 -269
-742 408
-427 228
-281 146
172 -86
-663 323
-460 217
-358 164
-268 118
5 -2
-432 179
65 -26
-701 270
-487 181
-433 155
-389 133
-357 118
-263 83
-436 132
-373 108
-357 98
-323 85
-294 73
-362 86
-328 73
-309 65
-336 66
-321 59
-320 55
-309 49
-313 46
-309 41
-304 37
-307 34
-301 29
-299 25
-303 22
-290 17
-286 14
-287 10
-301 7
-297 3
-292 0
-297 -3
-301 -7
-287 -10
-286 -14
-290 -17
-303 -22
-299 -25
-301 -29
-307 -34
-304 -37
-309 -41
-313 -46
-309 -49
-320 -55
-321 -59
-336 -66
-309 -65
-328 -73
-362 -86
-294 -73
-323 -85
-357 -98
-373 -108
-436 -132
-263 -83
-357 -118
-389 -133
-433 -155
-487 -181
-701 -270
65 26
-432 -179
5 2
-268 -118
-358 -164
-460 -217
-663 -323
172 86
-281 -146
-427 -228
-742 -408
476 269
-170 -99
-291 -174
-382 -235
-450 -285
-538 -350
-695 -464
-1166 -800
1116 786
-226 -163
-536 -397
-902 -686
-2022 -1578
4419 3536
791 649
304 255
76 66
-56 -50
-168 -153
-287 -266
-411 -391
-597 -582
-906 -906
-1765 -1809
2039 2141
2943 3168
3925 4331
1117 1263
683 792
478 569
345 420
236 295
116 148
-146 -191
1711 2307
428 593
285 405
227 331
173 260
142 219
98 155
60 98
-31 -51
680 1168
91 160
615 1118
166 311
112 216
75 150
11 23
606 1282
145 317
105 238
86 201
68 164
64 162
58 151
51 139
47 132
39 115
36 110
28 91
66 218
30 103
23 84
22 86
35 142
20 87
14 64
13 65
17 90
11 59
9 56
6 39
8 59
5 42
3 30
4 44
3 32
1 16
1 25
1 26
1 21
0 6
0 14
0 10
