0 0
0 -3
0 -9
2 -19
6 -30
11 -45
12 -40
19 -53
24 -59
36 -77
53 -100
83 -139
289 -432
51 -69
141 -172
478 -527
498 -498
587 -532
198 -162
-195 145
-196 130
-277 166
-90 48
-275 130
-184 76
-204 73
-173 52
-167 41
-167 33
-167 24
-159 15
-157 7
-156 0
-157 -7
-159 -15
-167 -24
-167 -33
-167 -41
-173 -52
-204 -73
-184 -76
-275 -130
-90 -48
-277 -166
-196 -130
-195 -145
198 162
587 532
498 498
478 527
141 172
51 69
289 432
83 139
53 100
36 77
24 59
19 53
12 40
11 45
6 30
2 19
0 9
0 3
