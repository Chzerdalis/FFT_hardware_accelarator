gen_input_real[0] = 32'sd0;
gen_input_real[16] = 32'sd32767;
gen_input_real[32] = -32'sd6738;
gen_input_real[48] = -32'sd24327;
gen_input_real[4] = 32'sd9756;
gen_input_real[20] = 32'sd15217;
gen_input_real[36] = -32'sd10062;
gen_input_real[52] = -32'sd7920;
gen_input_real[8] = 32'sd10717;
gen_input_real[24] = 32'sd3571;
gen_input_real[40] = -32'sd11792;
gen_input_real[56] = -32'sd1924;
gen_input_real[12] = 32'sd10901;
gen_input_real[28] = 32'sd958;
gen_input_real[44] = -32'sd7267;
gen_input_real[60] = -32'sd1439;
gen_input_real[1] = 32'sd2208;
gen_input_real[17] = 32'sd2554;
gen_input_real[33] = 32'sd2413;
gen_input_real[49] = -32'sd1936;
gen_input_real[5] = -32'sd4438;
gen_input_real[21] = -32'sd699;
gen_input_real[37] = 32'sd4139;
gen_input_real[53] = 32'sd4303;
gen_input_real[9] = -32'sd3791;
gen_input_real[25] = -32'sd6510;
gen_input_real[41] = 32'sd3481;
gen_input_real[57] = 32'sd4526;
gen_input_real[13] = -32'sd2133;
gen_input_real[29] = 32'sd594;
gen_input_real[45] = -32'sd783;
gen_input_real[61] = -32'sd3037;
gen_input_real[2] = 32'sd3037;
gen_input_real[18] = 32'sd783;
gen_input_real[34] = -32'sd594;
gen_input_real[50] = 32'sd2133;
gen_input_real[6] = -32'sd4526;
gen_input_real[22] = -32'sd3481;
gen_input_real[38] = 32'sd6510;
gen_input_real[54] = 32'sd3791;
gen_input_real[10] = -32'sd4303;
gen_input_real[26] = -32'sd4139;
gen_input_real[42] = 32'sd699;
gen_input_real[58] = 32'sd4438;
gen_input_real[14] = 32'sd1936;
gen_input_real[30] = -32'sd2413;
gen_input_real[46] = -32'sd2554;
gen_input_real[62] = -32'sd2208;
gen_input_real[3] = 32'sd1439;
gen_input_real[19] = 32'sd7267;
gen_input_real[35] = -32'sd958;
gen_input_real[51] = -32'sd10901;
gen_input_real[7] = 32'sd1924;
gen_input_real[23] = 32'sd11792;
gen_input_real[39] = -32'sd3571;
gen_input_real[55] = -32'sd10717;
gen_input_real[11] = 32'sd7920;
gen_input_real[27] = 32'sd10062;
gen_input_real[43] = -32'sd15217;
gen_input_real[59] = -32'sd9756;
gen_input_real[15] = 32'sd24327;
gen_input_real[31] = 32'sd6738;
gen_input_real[47] = -32'sd32767;
gen_input_real[63] = 32'sd0;
