0 0
1388 -6980
8723 -21060
30011 -44915
117582 -117582
-47253 31573
-44173 18297
-45531 9056
-41496 0
-45531 -9056
-44173 -18297
-47253 -31573
117582 117582
30011 44915
8723 21060
1388 6980
