w_real[0] = 9'h0FF; w_imag[0] = 9'h000;
w_real[1] = 9'h0FF; w_imag[1] = 9'h1FF;
w_real[2] = 9'h0FF; w_imag[2] = 9'h1FD;
w_real[3] = 9'h0FF; w_imag[3] = 9'h1FC;
w_real[4] = 9'h0FF; w_imag[4] = 9'h1FA;
w_real[5] = 9'h0FF; w_imag[5] = 9'h1F9;
w_real[6] = 9'h0FF; w_imag[6] = 9'h1F7;
w_real[7] = 9'h0FF; w_imag[7] = 9'h1F6;
w_real[8] = 9'h0FF; w_imag[8] = 9'h1F4;
w_real[9] = 9'h0FF; w_imag[9] = 9'h1F2;
w_real[10] = 9'h0FF; w_imag[10] = 9'h1F1;
w_real[11] = 9'h0FF; w_imag[11] = 9'h1EF;
w_real[12] = 9'h0FF; w_imag[12] = 9'h1EE;
w_real[13] = 9'h0FF; w_imag[13] = 9'h1EC;
w_real[14] = 9'h0FF; w_imag[14] = 9'h1EB;
w_real[15] = 9'h0FE; w_imag[15] = 9'h1E9;
w_real[16] = 9'h0FE; w_imag[16] = 9'h1E7;
w_real[17] = 9'h0FE; w_imag[17] = 9'h1E6;
w_real[18] = 9'h0FE; w_imag[18] = 9'h1E4;
w_real[19] = 9'h0FE; w_imag[19] = 9'h1E3;
w_real[20] = 9'h0FE; w_imag[20] = 9'h1E1;
w_real[21] = 9'h0FD; w_imag[21] = 9'h1E0;
w_real[22] = 9'h0FD; w_imag[22] = 9'h1DE;
w_real[23] = 9'h0FD; w_imag[23] = 9'h1DC;
w_real[24] = 9'h0FD; w_imag[24] = 9'h1DB;
w_real[25] = 9'h0FC; w_imag[25] = 9'h1D9;
w_real[26] = 9'h0FC; w_imag[26] = 9'h1D8;
w_real[27] = 9'h0FC; w_imag[27] = 9'h1D6;
w_real[28] = 9'h0FC; w_imag[28] = 9'h1D5;
w_real[29] = 9'h0FB; w_imag[29] = 9'h1D3;
w_real[30] = 9'h0FB; w_imag[30] = 9'h1D2;
w_real[31] = 9'h0FB; w_imag[31] = 9'h1D0;
w_real[32] = 9'h0FB; w_imag[32] = 9'h1CF;
w_real[33] = 9'h0FA; w_imag[33] = 9'h1CD;
w_real[34] = 9'h0FA; w_imag[34] = 9'h1CB;
w_real[35] = 9'h0FA; w_imag[35] = 9'h1CA;
w_real[36] = 9'h0F9; w_imag[36] = 9'h1C8;
w_real[37] = 9'h0F9; w_imag[37] = 9'h1C7;
w_real[38] = 9'h0F9; w_imag[38] = 9'h1C5;
w_real[39] = 9'h0F8; w_imag[39] = 9'h1C4;
w_real[40] = 9'h0F8; w_imag[40] = 9'h1C2;
w_real[41] = 9'h0F7; w_imag[41] = 9'h1C1;
w_real[42] = 9'h0F7; w_imag[42] = 9'h1BF;
w_real[43] = 9'h0F7; w_imag[43] = 9'h1BE;
w_real[44] = 9'h0F6; w_imag[44] = 9'h1BC;
w_real[45] = 9'h0F6; w_imag[45] = 9'h1BB;
w_real[46] = 9'h0F5; w_imag[46] = 9'h1B9;
w_real[47] = 9'h0F5; w_imag[47] = 9'h1B8;
w_real[48] = 9'h0F4; w_imag[48] = 9'h1B6;
w_real[49] = 9'h0F4; w_imag[49] = 9'h1B5;
w_real[50] = 9'h0F4; w_imag[50] = 9'h1B3;
w_real[51] = 9'h0F3; w_imag[51] = 9'h1B2;
w_real[52] = 9'h0F3; w_imag[52] = 9'h1B0;
w_real[53] = 9'h0F2; w_imag[53] = 9'h1AF;
w_real[54] = 9'h0F2; w_imag[54] = 9'h1AD;
w_real[55] = 9'h0F1; w_imag[55] = 9'h1AC;
w_real[56] = 9'h0F1; w_imag[56] = 9'h1AA;
w_real[57] = 9'h0F0; w_imag[57] = 9'h1A9;
w_real[58] = 9'h0EF; w_imag[58] = 9'h1A7;
w_real[59] = 9'h0EF; w_imag[59] = 9'h1A6;
w_real[60] = 9'h0EE; w_imag[60] = 9'h1A4;
w_real[61] = 9'h0EE; w_imag[61] = 9'h1A3;
w_real[62] = 9'h0ED; w_imag[62] = 9'h1A1;
w_real[63] = 9'h0ED; w_imag[63] = 9'h1A0;
w_real[64] = 9'h0EC; w_imag[64] = 9'h19F;
w_real[65] = 9'h0EB; w_imag[65] = 9'h19D;
w_real[66] = 9'h0EB; w_imag[66] = 9'h19C;
w_real[67] = 9'h0EA; w_imag[67] = 9'h19A;
w_real[68] = 9'h0EA; w_imag[68] = 9'h199;
w_real[69] = 9'h0E9; w_imag[69] = 9'h197;
w_real[70] = 9'h0E8; w_imag[70] = 9'h196;
w_real[71] = 9'h0E8; w_imag[71] = 9'h194;
w_real[72] = 9'h0E7; w_imag[72] = 9'h193;
w_real[73] = 9'h0E6; w_imag[73] = 9'h192;
w_real[74] = 9'h0E6; w_imag[74] = 9'h190;
w_real[75] = 9'h0E5; w_imag[75] = 9'h18F;
w_real[76] = 9'h0E4; w_imag[76] = 9'h18D;
w_real[77] = 9'h0E3; w_imag[77] = 9'h18C;
w_real[78] = 9'h0E3; w_imag[78] = 9'h18B;
w_real[79] = 9'h0E2; w_imag[79] = 9'h189;
w_real[80] = 9'h0E1; w_imag[80] = 9'h188;
w_real[81] = 9'h0E1; w_imag[81] = 9'h186;
w_real[82] = 9'h0E0; w_imag[82] = 9'h185;
w_real[83] = 9'h0DF; w_imag[83] = 9'h184;
w_real[84] = 9'h0DE; w_imag[84] = 9'h182;
w_real[85] = 9'h0DD; w_imag[85] = 9'h181;
w_real[86] = 9'h0DD; w_imag[86] = 9'h180;
w_real[87] = 9'h0DC; w_imag[87] = 9'h17E;
w_real[88] = 9'h0DB; w_imag[88] = 9'h17D;
w_real[89] = 9'h0DA; w_imag[89] = 9'h17C;
w_real[90] = 9'h0D9; w_imag[90] = 9'h17A;
w_real[91] = 9'h0D9; w_imag[91] = 9'h179;
w_real[92] = 9'h0D8; w_imag[92] = 9'h178;
w_real[93] = 9'h0D7; w_imag[93] = 9'h176;
w_real[94] = 9'h0D6; w_imag[94] = 9'h175;
w_real[95] = 9'h0D5; w_imag[95] = 9'h174;
w_real[96] = 9'h0D4; w_imag[96] = 9'h172;
w_real[97] = 9'h0D3; w_imag[97] = 9'h171;
w_real[98] = 9'h0D3; w_imag[98] = 9'h170;
w_real[99] = 9'h0D2; w_imag[99] = 9'h16E;
w_real[100] = 9'h0D1; w_imag[100] = 9'h16D;
w_real[101] = 9'h0D0; w_imag[101] = 9'h16C;
w_real[102] = 9'h0CF; w_imag[102] = 9'h16B;
w_real[103] = 9'h0CE; w_imag[103] = 9'h169;
w_real[104] = 9'h0CD; w_imag[104] = 9'h168;
w_real[105] = 9'h0CC; w_imag[105] = 9'h167;
w_real[106] = 9'h0CB; w_imag[106] = 9'h165;
w_real[107] = 9'h0CA; w_imag[107] = 9'h164;
w_real[108] = 9'h0C9; w_imag[108] = 9'h163;
w_real[109] = 9'h0C8; w_imag[109] = 9'h162;
w_real[110] = 9'h0C7; w_imag[110] = 9'h161;
w_real[111] = 9'h0C6; w_imag[111] = 9'h15F;
w_real[112] = 9'h0C5; w_imag[112] = 9'h15E;
w_real[113] = 9'h0C4; w_imag[113] = 9'h15D;
w_real[114] = 9'h0C3; w_imag[114] = 9'h15C;
w_real[115] = 9'h0C2; w_imag[115] = 9'h15A;
w_real[116] = 9'h0C1; w_imag[116] = 9'h159;
w_real[117] = 9'h0C0; w_imag[117] = 9'h158;
w_real[118] = 9'h0BF; w_imag[118] = 9'h157;
w_real[119] = 9'h0BE; w_imag[119] = 9'h156;
w_real[120] = 9'h0BD; w_imag[120] = 9'h155;
w_real[121] = 9'h0BC; w_imag[121] = 9'h153;
w_real[122] = 9'h0BB; w_imag[122] = 9'h152;
w_real[123] = 9'h0BA; w_imag[123] = 9'h151;
w_real[124] = 9'h0B9; w_imag[124] = 9'h150;
w_real[125] = 9'h0B8; w_imag[125] = 9'h14F;
w_real[126] = 9'h0B7; w_imag[126] = 9'h14E;
w_real[127] = 9'h0B6; w_imag[127] = 9'h14D;
w_real[128] = 9'h0B5; w_imag[128] = 9'h14B;
w_real[129] = 9'h0B3; w_imag[129] = 9'h14A;
w_real[130] = 9'h0B2; w_imag[130] = 9'h149;
w_real[131] = 9'h0B1; w_imag[131] = 9'h148;
w_real[132] = 9'h0B0; w_imag[132] = 9'h147;
w_real[133] = 9'h0AF; w_imag[133] = 9'h146;
w_real[134] = 9'h0AE; w_imag[134] = 9'h145;
w_real[135] = 9'h0AD; w_imag[135] = 9'h144;
w_real[136] = 9'h0AB; w_imag[136] = 9'h143;
w_real[137] = 9'h0AA; w_imag[137] = 9'h142;
w_real[138] = 9'h0A9; w_imag[138] = 9'h141;
w_real[139] = 9'h0A8; w_imag[139] = 9'h140;
w_real[140] = 9'h0A7; w_imag[140] = 9'h13F;
w_real[141] = 9'h0A6; w_imag[141] = 9'h13E;
w_real[142] = 9'h0A4; w_imag[142] = 9'h13D;
w_real[143] = 9'h0A3; w_imag[143] = 9'h13C;
w_real[144] = 9'h0A2; w_imag[144] = 9'h13B;
w_real[145] = 9'h0A1; w_imag[145] = 9'h13A;
w_real[146] = 9'h09F; w_imag[146] = 9'h139;
w_real[147] = 9'h09E; w_imag[147] = 9'h138;
w_real[148] = 9'h09D; w_imag[148] = 9'h137;
w_real[149] = 9'h09C; w_imag[149] = 9'h136;
w_real[150] = 9'h09B; w_imag[150] = 9'h135;
w_real[151] = 9'h099; w_imag[151] = 9'h134;
w_real[152] = 9'h098; w_imag[152] = 9'h133;
w_real[153] = 9'h097; w_imag[153] = 9'h132;
w_real[154] = 9'h095; w_imag[154] = 9'h131;
w_real[155] = 9'h094; w_imag[155] = 9'h130;
w_real[156] = 9'h093; w_imag[156] = 9'h12F;
w_real[157] = 9'h092; w_imag[157] = 9'h12E;
w_real[158] = 9'h090; w_imag[158] = 9'h12D;
w_real[159] = 9'h08F; w_imag[159] = 9'h12D;
w_real[160] = 9'h08E; w_imag[160] = 9'h12C;
w_real[161] = 9'h08C; w_imag[161] = 9'h12B;
w_real[162] = 9'h08B; w_imag[162] = 9'h12A;
w_real[163] = 9'h08A; w_imag[163] = 9'h129;
w_real[164] = 9'h088; w_imag[164] = 9'h128;
w_real[165] = 9'h087; w_imag[165] = 9'h127;
w_real[166] = 9'h086; w_imag[166] = 9'h127;
w_real[167] = 9'h084; w_imag[167] = 9'h126;
w_real[168] = 9'h083; w_imag[168] = 9'h125;
w_real[169] = 9'h082; w_imag[169] = 9'h124;
w_real[170] = 9'h080; w_imag[170] = 9'h123;
w_real[171] = 9'h07F; w_imag[171] = 9'h123;
w_real[172] = 9'h07E; w_imag[172] = 9'h122;
w_real[173] = 9'h07C; w_imag[173] = 9'h121;
w_real[174] = 9'h07B; w_imag[174] = 9'h120;
w_real[175] = 9'h07A; w_imag[175] = 9'h11F;
w_real[176] = 9'h078; w_imag[176] = 9'h11F;
w_real[177] = 9'h077; w_imag[177] = 9'h11E;
w_real[178] = 9'h075; w_imag[178] = 9'h11D;
w_real[179] = 9'h074; w_imag[179] = 9'h11D;
w_real[180] = 9'h073; w_imag[180] = 9'h11C;
w_real[181] = 9'h071; w_imag[181] = 9'h11B;
w_real[182] = 9'h070; w_imag[182] = 9'h11A;
w_real[183] = 9'h06E; w_imag[183] = 9'h11A;
w_real[184] = 9'h06D; w_imag[184] = 9'h119;
w_real[185] = 9'h06C; w_imag[185] = 9'h118;
w_real[186] = 9'h06A; w_imag[186] = 9'h118;
w_real[187] = 9'h069; w_imag[187] = 9'h117;
w_real[188] = 9'h067; w_imag[188] = 9'h116;
w_real[189] = 9'h066; w_imag[189] = 9'h116;
w_real[190] = 9'h064; w_imag[190] = 9'h115;
w_real[191] = 9'h063; w_imag[191] = 9'h115;
w_real[192] = 9'h061; w_imag[192] = 9'h114;
w_real[193] = 9'h060; w_imag[193] = 9'h113;
w_real[194] = 9'h05F; w_imag[194] = 9'h113;
w_real[195] = 9'h05D; w_imag[195] = 9'h112;
w_real[196] = 9'h05C; w_imag[196] = 9'h112;
w_real[197] = 9'h05A; w_imag[197] = 9'h111;
w_real[198] = 9'h059; w_imag[198] = 9'h111;
w_real[199] = 9'h057; w_imag[199] = 9'h110;
w_real[200] = 9'h056; w_imag[200] = 9'h10F;
w_real[201] = 9'h054; w_imag[201] = 9'h10F;
w_real[202] = 9'h053; w_imag[202] = 9'h10E;
w_real[203] = 9'h051; w_imag[203] = 9'h10E;
w_real[204] = 9'h050; w_imag[204] = 9'h10D;
w_real[205] = 9'h04E; w_imag[205] = 9'h10D;
w_real[206] = 9'h04D; w_imag[206] = 9'h10C;
w_real[207] = 9'h04B; w_imag[207] = 9'h10C;
w_real[208] = 9'h04A; w_imag[208] = 9'h10C;
w_real[209] = 9'h048; w_imag[209] = 9'h10B;
w_real[210] = 9'h047; w_imag[210] = 9'h10B;
w_real[211] = 9'h045; w_imag[211] = 9'h10A;
w_real[212] = 9'h044; w_imag[212] = 9'h10A;
w_real[213] = 9'h042; w_imag[213] = 9'h109;
w_real[214] = 9'h041; w_imag[214] = 9'h109;
w_real[215] = 9'h03F; w_imag[215] = 9'h109;
w_real[216] = 9'h03E; w_imag[216] = 9'h108;
w_real[217] = 9'h03C; w_imag[217] = 9'h108;
w_real[218] = 9'h03B; w_imag[218] = 9'h107;
w_real[219] = 9'h039; w_imag[219] = 9'h107;
w_real[220] = 9'h038; w_imag[220] = 9'h107;
w_real[221] = 9'h036; w_imag[221] = 9'h106;
w_real[222] = 9'h035; w_imag[222] = 9'h106;
w_real[223] = 9'h033; w_imag[223] = 9'h106;
w_real[224] = 9'h031; w_imag[224] = 9'h105;
w_real[225] = 9'h030; w_imag[225] = 9'h105;
w_real[226] = 9'h02E; w_imag[226] = 9'h105;
w_real[227] = 9'h02D; w_imag[227] = 9'h105;
w_real[228] = 9'h02B; w_imag[228] = 9'h104;
w_real[229] = 9'h02A; w_imag[229] = 9'h104;
w_real[230] = 9'h028; w_imag[230] = 9'h104;
w_real[231] = 9'h027; w_imag[231] = 9'h104;
w_real[232] = 9'h025; w_imag[232] = 9'h103;
w_real[233] = 9'h024; w_imag[233] = 9'h103;
w_real[234] = 9'h022; w_imag[234] = 9'h103;
w_real[235] = 9'h020; w_imag[235] = 9'h103;
w_real[236] = 9'h01F; w_imag[236] = 9'h102;
w_real[237] = 9'h01D; w_imag[237] = 9'h102;
w_real[238] = 9'h01C; w_imag[238] = 9'h102;
w_real[239] = 9'h01A; w_imag[239] = 9'h102;
w_real[240] = 9'h019; w_imag[240] = 9'h102;
w_real[241] = 9'h017; w_imag[241] = 9'h102;
w_real[242] = 9'h015; w_imag[242] = 9'h101;
w_real[243] = 9'h014; w_imag[243] = 9'h101;
w_real[244] = 9'h012; w_imag[244] = 9'h101;
w_real[245] = 9'h011; w_imag[245] = 9'h101;
w_real[246] = 9'h00F; w_imag[246] = 9'h101;
w_real[247] = 9'h00E; w_imag[247] = 9'h101;
w_real[248] = 9'h00C; w_imag[248] = 9'h101;
w_real[249] = 9'h00A; w_imag[249] = 9'h101;
w_real[250] = 9'h009; w_imag[250] = 9'h101;
w_real[251] = 9'h007; w_imag[251] = 9'h101;
w_real[252] = 9'h006; w_imag[252] = 9'h101;
w_real[253] = 9'h004; w_imag[253] = 9'h101;
w_real[254] = 9'h003; w_imag[254] = 9'h101;
w_real[255] = 9'h001; w_imag[255] = 9'h101;
w_real[256] = 9'h000; w_imag[256] = 9'h100;
w_real[257] = 9'h1FF; w_imag[257] = 9'h101;
w_real[258] = 9'h1FD; w_imag[258] = 9'h101;
w_real[259] = 9'h1FC; w_imag[259] = 9'h101;
w_real[260] = 9'h1FA; w_imag[260] = 9'h101;
w_real[261] = 9'h1F9; w_imag[261] = 9'h101;
w_real[262] = 9'h1F7; w_imag[262] = 9'h101;
w_real[263] = 9'h1F6; w_imag[263] = 9'h101;
w_real[264] = 9'h1F4; w_imag[264] = 9'h101;
w_real[265] = 9'h1F2; w_imag[265] = 9'h101;
w_real[266] = 9'h1F1; w_imag[266] = 9'h101;
w_real[267] = 9'h1EF; w_imag[267] = 9'h101;
w_real[268] = 9'h1EE; w_imag[268] = 9'h101;
w_real[269] = 9'h1EC; w_imag[269] = 9'h101;
w_real[270] = 9'h1EB; w_imag[270] = 9'h101;
w_real[271] = 9'h1E9; w_imag[271] = 9'h102;
w_real[272] = 9'h1E7; w_imag[272] = 9'h102;
w_real[273] = 9'h1E6; w_imag[273] = 9'h102;
w_real[274] = 9'h1E4; w_imag[274] = 9'h102;
w_real[275] = 9'h1E3; w_imag[275] = 9'h102;
w_real[276] = 9'h1E1; w_imag[276] = 9'h102;
w_real[277] = 9'h1E0; w_imag[277] = 9'h103;
w_real[278] = 9'h1DE; w_imag[278] = 9'h103;
w_real[279] = 9'h1DC; w_imag[279] = 9'h103;
w_real[280] = 9'h1DB; w_imag[280] = 9'h103;
w_real[281] = 9'h1D9; w_imag[281] = 9'h104;
w_real[282] = 9'h1D8; w_imag[282] = 9'h104;
w_real[283] = 9'h1D6; w_imag[283] = 9'h104;
w_real[284] = 9'h1D5; w_imag[284] = 9'h104;
w_real[285] = 9'h1D3; w_imag[285] = 9'h105;
w_real[286] = 9'h1D2; w_imag[286] = 9'h105;
w_real[287] = 9'h1D0; w_imag[287] = 9'h105;
w_real[288] = 9'h1CF; w_imag[288] = 9'h105;
w_real[289] = 9'h1CD; w_imag[289] = 9'h106;
w_real[290] = 9'h1CB; w_imag[290] = 9'h106;
w_real[291] = 9'h1CA; w_imag[291] = 9'h106;
w_real[292] = 9'h1C8; w_imag[292] = 9'h107;
w_real[293] = 9'h1C7; w_imag[293] = 9'h107;
w_real[294] = 9'h1C5; w_imag[294] = 9'h107;
w_real[295] = 9'h1C4; w_imag[295] = 9'h108;
w_real[296] = 9'h1C2; w_imag[296] = 9'h108;
w_real[297] = 9'h1C1; w_imag[297] = 9'h109;
w_real[298] = 9'h1BF; w_imag[298] = 9'h109;
w_real[299] = 9'h1BE; w_imag[299] = 9'h109;
w_real[300] = 9'h1BC; w_imag[300] = 9'h10A;
w_real[301] = 9'h1BB; w_imag[301] = 9'h10A;
w_real[302] = 9'h1B9; w_imag[302] = 9'h10B;
w_real[303] = 9'h1B8; w_imag[303] = 9'h10B;
w_real[304] = 9'h1B6; w_imag[304] = 9'h10C;
w_real[305] = 9'h1B5; w_imag[305] = 9'h10C;
w_real[306] = 9'h1B3; w_imag[306] = 9'h10C;
w_real[307] = 9'h1B2; w_imag[307] = 9'h10D;
w_real[308] = 9'h1B0; w_imag[308] = 9'h10D;
w_real[309] = 9'h1AF; w_imag[309] = 9'h10E;
w_real[310] = 9'h1AD; w_imag[310] = 9'h10E;
w_real[311] = 9'h1AC; w_imag[311] = 9'h10F;
w_real[312] = 9'h1AA; w_imag[312] = 9'h10F;
w_real[313] = 9'h1A9; w_imag[313] = 9'h110;
w_real[314] = 9'h1A7; w_imag[314] = 9'h111;
w_real[315] = 9'h1A6; w_imag[315] = 9'h111;
w_real[316] = 9'h1A4; w_imag[316] = 9'h112;
w_real[317] = 9'h1A3; w_imag[317] = 9'h112;
w_real[318] = 9'h1A1; w_imag[318] = 9'h113;
w_real[319] = 9'h1A0; w_imag[319] = 9'h113;
w_real[320] = 9'h19F; w_imag[320] = 9'h114;
w_real[321] = 9'h19D; w_imag[321] = 9'h115;
w_real[322] = 9'h19C; w_imag[322] = 9'h115;
w_real[323] = 9'h19A; w_imag[323] = 9'h116;
w_real[324] = 9'h199; w_imag[324] = 9'h116;
w_real[325] = 9'h197; w_imag[325] = 9'h117;
w_real[326] = 9'h196; w_imag[326] = 9'h118;
w_real[327] = 9'h194; w_imag[327] = 9'h118;
w_real[328] = 9'h193; w_imag[328] = 9'h119;
w_real[329] = 9'h192; w_imag[329] = 9'h11A;
w_real[330] = 9'h190; w_imag[330] = 9'h11A;
w_real[331] = 9'h18F; w_imag[331] = 9'h11B;
w_real[332] = 9'h18D; w_imag[332] = 9'h11C;
w_real[333] = 9'h18C; w_imag[333] = 9'h11D;
w_real[334] = 9'h18B; w_imag[334] = 9'h11D;
w_real[335] = 9'h189; w_imag[335] = 9'h11E;
w_real[336] = 9'h188; w_imag[336] = 9'h11F;
w_real[337] = 9'h186; w_imag[337] = 9'h11F;
w_real[338] = 9'h185; w_imag[338] = 9'h120;
w_real[339] = 9'h184; w_imag[339] = 9'h121;
w_real[340] = 9'h182; w_imag[340] = 9'h122;
w_real[341] = 9'h181; w_imag[341] = 9'h123;
w_real[342] = 9'h180; w_imag[342] = 9'h123;
w_real[343] = 9'h17E; w_imag[343] = 9'h124;
w_real[344] = 9'h17D; w_imag[344] = 9'h125;
w_real[345] = 9'h17C; w_imag[345] = 9'h126;
w_real[346] = 9'h17A; w_imag[346] = 9'h127;
w_real[347] = 9'h179; w_imag[347] = 9'h127;
w_real[348] = 9'h178; w_imag[348] = 9'h128;
w_real[349] = 9'h176; w_imag[349] = 9'h129;
w_real[350] = 9'h175; w_imag[350] = 9'h12A;
w_real[351] = 9'h174; w_imag[351] = 9'h12B;
w_real[352] = 9'h172; w_imag[352] = 9'h12C;
w_real[353] = 9'h171; w_imag[353] = 9'h12D;
w_real[354] = 9'h170; w_imag[354] = 9'h12D;
w_real[355] = 9'h16E; w_imag[355] = 9'h12E;
w_real[356] = 9'h16D; w_imag[356] = 9'h12F;
w_real[357] = 9'h16C; w_imag[357] = 9'h130;
w_real[358] = 9'h16B; w_imag[358] = 9'h131;
w_real[359] = 9'h169; w_imag[359] = 9'h132;
w_real[360] = 9'h168; w_imag[360] = 9'h133;
w_real[361] = 9'h167; w_imag[361] = 9'h134;
w_real[362] = 9'h165; w_imag[362] = 9'h135;
w_real[363] = 9'h164; w_imag[363] = 9'h136;
w_real[364] = 9'h163; w_imag[364] = 9'h137;
w_real[365] = 9'h162; w_imag[365] = 9'h138;
w_real[366] = 9'h161; w_imag[366] = 9'h139;
w_real[367] = 9'h15F; w_imag[367] = 9'h13A;
w_real[368] = 9'h15E; w_imag[368] = 9'h13B;
w_real[369] = 9'h15D; w_imag[369] = 9'h13C;
w_real[370] = 9'h15C; w_imag[370] = 9'h13D;
w_real[371] = 9'h15A; w_imag[371] = 9'h13E;
w_real[372] = 9'h159; w_imag[372] = 9'h13F;
w_real[373] = 9'h158; w_imag[373] = 9'h140;
w_real[374] = 9'h157; w_imag[374] = 9'h141;
w_real[375] = 9'h156; w_imag[375] = 9'h142;
w_real[376] = 9'h155; w_imag[376] = 9'h143;
w_real[377] = 9'h153; w_imag[377] = 9'h144;
w_real[378] = 9'h152; w_imag[378] = 9'h145;
w_real[379] = 9'h151; w_imag[379] = 9'h146;
w_real[380] = 9'h150; w_imag[380] = 9'h147;
w_real[381] = 9'h14F; w_imag[381] = 9'h148;
w_real[382] = 9'h14E; w_imag[382] = 9'h149;
w_real[383] = 9'h14D; w_imag[383] = 9'h14A;
w_real[384] = 9'h14B; w_imag[384] = 9'h14B;
w_real[385] = 9'h14A; w_imag[385] = 9'h14D;
w_real[386] = 9'h149; w_imag[386] = 9'h14E;
w_real[387] = 9'h148; w_imag[387] = 9'h14F;
w_real[388] = 9'h147; w_imag[388] = 9'h150;
w_real[389] = 9'h146; w_imag[389] = 9'h151;
w_real[390] = 9'h145; w_imag[390] = 9'h152;
w_real[391] = 9'h144; w_imag[391] = 9'h153;
w_real[392] = 9'h143; w_imag[392] = 9'h155;
w_real[393] = 9'h142; w_imag[393] = 9'h156;
w_real[394] = 9'h141; w_imag[394] = 9'h157;
w_real[395] = 9'h140; w_imag[395] = 9'h158;
w_real[396] = 9'h13F; w_imag[396] = 9'h159;
w_real[397] = 9'h13E; w_imag[397] = 9'h15A;
w_real[398] = 9'h13D; w_imag[398] = 9'h15C;
w_real[399] = 9'h13C; w_imag[399] = 9'h15D;
w_real[400] = 9'h13B; w_imag[400] = 9'h15E;
w_real[401] = 9'h13A; w_imag[401] = 9'h15F;
w_real[402] = 9'h139; w_imag[402] = 9'h161;
w_real[403] = 9'h138; w_imag[403] = 9'h162;
w_real[404] = 9'h137; w_imag[404] = 9'h163;
w_real[405] = 9'h136; w_imag[405] = 9'h164;
w_real[406] = 9'h135; w_imag[406] = 9'h165;
w_real[407] = 9'h134; w_imag[407] = 9'h167;
w_real[408] = 9'h133; w_imag[408] = 9'h168;
w_real[409] = 9'h132; w_imag[409] = 9'h169;
w_real[410] = 9'h131; w_imag[410] = 9'h16B;
w_real[411] = 9'h130; w_imag[411] = 9'h16C;
w_real[412] = 9'h12F; w_imag[412] = 9'h16D;
w_real[413] = 9'h12E; w_imag[413] = 9'h16E;
w_real[414] = 9'h12D; w_imag[414] = 9'h170;
w_real[415] = 9'h12D; w_imag[415] = 9'h171;
w_real[416] = 9'h12C; w_imag[416] = 9'h172;
w_real[417] = 9'h12B; w_imag[417] = 9'h174;
w_real[418] = 9'h12A; w_imag[418] = 9'h175;
w_real[419] = 9'h129; w_imag[419] = 9'h176;
w_real[420] = 9'h128; w_imag[420] = 9'h178;
w_real[421] = 9'h127; w_imag[421] = 9'h179;
w_real[422] = 9'h127; w_imag[422] = 9'h17A;
w_real[423] = 9'h126; w_imag[423] = 9'h17C;
w_real[424] = 9'h125; w_imag[424] = 9'h17D;
w_real[425] = 9'h124; w_imag[425] = 9'h17E;
w_real[426] = 9'h123; w_imag[426] = 9'h180;
w_real[427] = 9'h123; w_imag[427] = 9'h181;
w_real[428] = 9'h122; w_imag[428] = 9'h182;
w_real[429] = 9'h121; w_imag[429] = 9'h184;
w_real[430] = 9'h120; w_imag[430] = 9'h185;
w_real[431] = 9'h11F; w_imag[431] = 9'h186;
w_real[432] = 9'h11F; w_imag[432] = 9'h188;
w_real[433] = 9'h11E; w_imag[433] = 9'h189;
w_real[434] = 9'h11D; w_imag[434] = 9'h18B;
w_real[435] = 9'h11D; w_imag[435] = 9'h18C;
w_real[436] = 9'h11C; w_imag[436] = 9'h18D;
w_real[437] = 9'h11B; w_imag[437] = 9'h18F;
w_real[438] = 9'h11A; w_imag[438] = 9'h190;
w_real[439] = 9'h11A; w_imag[439] = 9'h192;
w_real[440] = 9'h119; w_imag[440] = 9'h193;
w_real[441] = 9'h118; w_imag[441] = 9'h194;
w_real[442] = 9'h118; w_imag[442] = 9'h196;
w_real[443] = 9'h117; w_imag[443] = 9'h197;
w_real[444] = 9'h116; w_imag[444] = 9'h199;
w_real[445] = 9'h116; w_imag[445] = 9'h19A;
w_real[446] = 9'h115; w_imag[446] = 9'h19C;
w_real[447] = 9'h115; w_imag[447] = 9'h19D;
w_real[448] = 9'h114; w_imag[448] = 9'h19F;
w_real[449] = 9'h113; w_imag[449] = 9'h1A0;
w_real[450] = 9'h113; w_imag[450] = 9'h1A1;
w_real[451] = 9'h112; w_imag[451] = 9'h1A3;
w_real[452] = 9'h112; w_imag[452] = 9'h1A4;
w_real[453] = 9'h111; w_imag[453] = 9'h1A6;
w_real[454] = 9'h111; w_imag[454] = 9'h1A7;
w_real[455] = 9'h110; w_imag[455] = 9'h1A9;
w_real[456] = 9'h10F; w_imag[456] = 9'h1AA;
w_real[457] = 9'h10F; w_imag[457] = 9'h1AC;
w_real[458] = 9'h10E; w_imag[458] = 9'h1AD;
w_real[459] = 9'h10E; w_imag[459] = 9'h1AF;
w_real[460] = 9'h10D; w_imag[460] = 9'h1B0;
w_real[461] = 9'h10D; w_imag[461] = 9'h1B2;
w_real[462] = 9'h10C; w_imag[462] = 9'h1B3;
w_real[463] = 9'h10C; w_imag[463] = 9'h1B5;
w_real[464] = 9'h10C; w_imag[464] = 9'h1B6;
w_real[465] = 9'h10B; w_imag[465] = 9'h1B8;
w_real[466] = 9'h10B; w_imag[466] = 9'h1B9;
w_real[467] = 9'h10A; w_imag[467] = 9'h1BB;
w_real[468] = 9'h10A; w_imag[468] = 9'h1BC;
w_real[469] = 9'h109; w_imag[469] = 9'h1BE;
w_real[470] = 9'h109; w_imag[470] = 9'h1BF;
w_real[471] = 9'h109; w_imag[471] = 9'h1C1;
w_real[472] = 9'h108; w_imag[472] = 9'h1C2;
w_real[473] = 9'h108; w_imag[473] = 9'h1C4;
w_real[474] = 9'h107; w_imag[474] = 9'h1C5;
w_real[475] = 9'h107; w_imag[475] = 9'h1C7;
w_real[476] = 9'h107; w_imag[476] = 9'h1C8;
w_real[477] = 9'h106; w_imag[477] = 9'h1CA;
w_real[478] = 9'h106; w_imag[478] = 9'h1CB;
w_real[479] = 9'h106; w_imag[479] = 9'h1CD;
w_real[480] = 9'h105; w_imag[480] = 9'h1CF;
w_real[481] = 9'h105; w_imag[481] = 9'h1D0;
w_real[482] = 9'h105; w_imag[482] = 9'h1D2;
w_real[483] = 9'h105; w_imag[483] = 9'h1D3;
w_real[484] = 9'h104; w_imag[484] = 9'h1D5;
w_real[485] = 9'h104; w_imag[485] = 9'h1D6;
w_real[486] = 9'h104; w_imag[486] = 9'h1D8;
w_real[487] = 9'h104; w_imag[487] = 9'h1D9;
w_real[488] = 9'h103; w_imag[488] = 9'h1DB;
w_real[489] = 9'h103; w_imag[489] = 9'h1DC;
w_real[490] = 9'h103; w_imag[490] = 9'h1DE;
w_real[491] = 9'h103; w_imag[491] = 9'h1E0;
w_real[492] = 9'h102; w_imag[492] = 9'h1E1;
w_real[493] = 9'h102; w_imag[493] = 9'h1E3;
w_real[494] = 9'h102; w_imag[494] = 9'h1E4;
w_real[495] = 9'h102; w_imag[495] = 9'h1E6;
w_real[496] = 9'h102; w_imag[496] = 9'h1E7;
w_real[497] = 9'h102; w_imag[497] = 9'h1E9;
w_real[498] = 9'h101; w_imag[498] = 9'h1EB;
w_real[499] = 9'h101; w_imag[499] = 9'h1EC;
w_real[500] = 9'h101; w_imag[500] = 9'h1EE;
w_real[501] = 9'h101; w_imag[501] = 9'h1EF;
w_real[502] = 9'h101; w_imag[502] = 9'h1F1;
w_real[503] = 9'h101; w_imag[503] = 9'h1F2;
w_real[504] = 9'h101; w_imag[504] = 9'h1F4;
w_real[505] = 9'h101; w_imag[505] = 9'h1F6;
w_real[506] = 9'h101; w_imag[506] = 9'h1F7;
w_real[507] = 9'h101; w_imag[507] = 9'h1F9;
w_real[508] = 9'h101; w_imag[508] = 9'h1FA;
w_real[509] = 9'h101; w_imag[509] = 9'h1FC;
w_real[510] = 9'h101; w_imag[510] = 9'h1FD;
w_real[511] = 9'h101; w_imag[511] = 9'h1FF;
w_real[512] = 9'h100; w_imag[512] = 9'h000;
w_real[513] = 9'h101; w_imag[513] = 9'h001;
w_real[514] = 9'h101; w_imag[514] = 9'h003;
w_real[515] = 9'h101; w_imag[515] = 9'h004;
w_real[516] = 9'h101; w_imag[516] = 9'h006;
w_real[517] = 9'h101; w_imag[517] = 9'h007;
w_real[518] = 9'h101; w_imag[518] = 9'h009;
w_real[519] = 9'h101; w_imag[519] = 9'h00A;
w_real[520] = 9'h101; w_imag[520] = 9'h00C;
w_real[521] = 9'h101; w_imag[521] = 9'h00E;
w_real[522] = 9'h101; w_imag[522] = 9'h00F;
w_real[523] = 9'h101; w_imag[523] = 9'h011;
w_real[524] = 9'h101; w_imag[524] = 9'h012;
w_real[525] = 9'h101; w_imag[525] = 9'h014;
w_real[526] = 9'h101; w_imag[526] = 9'h015;
w_real[527] = 9'h102; w_imag[527] = 9'h017;
w_real[528] = 9'h102; w_imag[528] = 9'h019;
w_real[529] = 9'h102; w_imag[529] = 9'h01A;
w_real[530] = 9'h102; w_imag[530] = 9'h01C;
w_real[531] = 9'h102; w_imag[531] = 9'h01D;
w_real[532] = 9'h102; w_imag[532] = 9'h01F;
w_real[533] = 9'h103; w_imag[533] = 9'h020;
w_real[534] = 9'h103; w_imag[534] = 9'h022;
w_real[535] = 9'h103; w_imag[535] = 9'h024;
w_real[536] = 9'h103; w_imag[536] = 9'h025;
w_real[537] = 9'h104; w_imag[537] = 9'h027;
w_real[538] = 9'h104; w_imag[538] = 9'h028;
w_real[539] = 9'h104; w_imag[539] = 9'h02A;
w_real[540] = 9'h104; w_imag[540] = 9'h02B;
w_real[541] = 9'h105; w_imag[541] = 9'h02D;
w_real[542] = 9'h105; w_imag[542] = 9'h02E;
w_real[543] = 9'h105; w_imag[543] = 9'h030;
w_real[544] = 9'h105; w_imag[544] = 9'h031;
w_real[545] = 9'h106; w_imag[545] = 9'h033;
w_real[546] = 9'h106; w_imag[546] = 9'h035;
w_real[547] = 9'h106; w_imag[547] = 9'h036;
w_real[548] = 9'h107; w_imag[548] = 9'h038;
w_real[549] = 9'h107; w_imag[549] = 9'h039;
w_real[550] = 9'h107; w_imag[550] = 9'h03B;
w_real[551] = 9'h108; w_imag[551] = 9'h03C;
w_real[552] = 9'h108; w_imag[552] = 9'h03E;
w_real[553] = 9'h109; w_imag[553] = 9'h03F;
w_real[554] = 9'h109; w_imag[554] = 9'h041;
w_real[555] = 9'h109; w_imag[555] = 9'h042;
w_real[556] = 9'h10A; w_imag[556] = 9'h044;
w_real[557] = 9'h10A; w_imag[557] = 9'h045;
w_real[558] = 9'h10B; w_imag[558] = 9'h047;
w_real[559] = 9'h10B; w_imag[559] = 9'h048;
w_real[560] = 9'h10C; w_imag[560] = 9'h04A;
w_real[561] = 9'h10C; w_imag[561] = 9'h04B;
w_real[562] = 9'h10C; w_imag[562] = 9'h04D;
w_real[563] = 9'h10D; w_imag[563] = 9'h04E;
w_real[564] = 9'h10D; w_imag[564] = 9'h050;
w_real[565] = 9'h10E; w_imag[565] = 9'h051;
w_real[566] = 9'h10E; w_imag[566] = 9'h053;
w_real[567] = 9'h10F; w_imag[567] = 9'h054;
w_real[568] = 9'h10F; w_imag[568] = 9'h056;
w_real[569] = 9'h110; w_imag[569] = 9'h057;
w_real[570] = 9'h111; w_imag[570] = 9'h059;
w_real[571] = 9'h111; w_imag[571] = 9'h05A;
w_real[572] = 9'h112; w_imag[572] = 9'h05C;
w_real[573] = 9'h112; w_imag[573] = 9'h05D;
w_real[574] = 9'h113; w_imag[574] = 9'h05F;
w_real[575] = 9'h113; w_imag[575] = 9'h060;
w_real[576] = 9'h114; w_imag[576] = 9'h061;
w_real[577] = 9'h115; w_imag[577] = 9'h063;
w_real[578] = 9'h115; w_imag[578] = 9'h064;
w_real[579] = 9'h116; w_imag[579] = 9'h066;
w_real[580] = 9'h116; w_imag[580] = 9'h067;
w_real[581] = 9'h117; w_imag[581] = 9'h069;
w_real[582] = 9'h118; w_imag[582] = 9'h06A;
w_real[583] = 9'h118; w_imag[583] = 9'h06C;
w_real[584] = 9'h119; w_imag[584] = 9'h06D;
w_real[585] = 9'h11A; w_imag[585] = 9'h06E;
w_real[586] = 9'h11A; w_imag[586] = 9'h070;
w_real[587] = 9'h11B; w_imag[587] = 9'h071;
w_real[588] = 9'h11C; w_imag[588] = 9'h073;
w_real[589] = 9'h11D; w_imag[589] = 9'h074;
w_real[590] = 9'h11D; w_imag[590] = 9'h075;
w_real[591] = 9'h11E; w_imag[591] = 9'h077;
w_real[592] = 9'h11F; w_imag[592] = 9'h078;
w_real[593] = 9'h11F; w_imag[593] = 9'h07A;
w_real[594] = 9'h120; w_imag[594] = 9'h07B;
w_real[595] = 9'h121; w_imag[595] = 9'h07C;
w_real[596] = 9'h122; w_imag[596] = 9'h07E;
w_real[597] = 9'h123; w_imag[597] = 9'h07F;
w_real[598] = 9'h123; w_imag[598] = 9'h080;
w_real[599] = 9'h124; w_imag[599] = 9'h082;
w_real[600] = 9'h125; w_imag[600] = 9'h083;
w_real[601] = 9'h126; w_imag[601] = 9'h084;
w_real[602] = 9'h127; w_imag[602] = 9'h086;
w_real[603] = 9'h127; w_imag[603] = 9'h087;
w_real[604] = 9'h128; w_imag[604] = 9'h088;
w_real[605] = 9'h129; w_imag[605] = 9'h08A;
w_real[606] = 9'h12A; w_imag[606] = 9'h08B;
w_real[607] = 9'h12B; w_imag[607] = 9'h08C;
w_real[608] = 9'h12C; w_imag[608] = 9'h08E;
w_real[609] = 9'h12D; w_imag[609] = 9'h08F;
w_real[610] = 9'h12D; w_imag[610] = 9'h090;
w_real[611] = 9'h12E; w_imag[611] = 9'h092;
w_real[612] = 9'h12F; w_imag[612] = 9'h093;
w_real[613] = 9'h130; w_imag[613] = 9'h094;
w_real[614] = 9'h131; w_imag[614] = 9'h095;
w_real[615] = 9'h132; w_imag[615] = 9'h097;
w_real[616] = 9'h133; w_imag[616] = 9'h098;
w_real[617] = 9'h134; w_imag[617] = 9'h099;
w_real[618] = 9'h135; w_imag[618] = 9'h09B;
w_real[619] = 9'h136; w_imag[619] = 9'h09C;
w_real[620] = 9'h137; w_imag[620] = 9'h09D;
w_real[621] = 9'h138; w_imag[621] = 9'h09E;
w_real[622] = 9'h139; w_imag[622] = 9'h09F;
w_real[623] = 9'h13A; w_imag[623] = 9'h0A1;
w_real[624] = 9'h13B; w_imag[624] = 9'h0A2;
w_real[625] = 9'h13C; w_imag[625] = 9'h0A3;
w_real[626] = 9'h13D; w_imag[626] = 9'h0A4;
w_real[627] = 9'h13E; w_imag[627] = 9'h0A6;
w_real[628] = 9'h13F; w_imag[628] = 9'h0A7;
w_real[629] = 9'h140; w_imag[629] = 9'h0A8;
w_real[630] = 9'h141; w_imag[630] = 9'h0A9;
w_real[631] = 9'h142; w_imag[631] = 9'h0AA;
w_real[632] = 9'h143; w_imag[632] = 9'h0AB;
w_real[633] = 9'h144; w_imag[633] = 9'h0AD;
w_real[634] = 9'h145; w_imag[634] = 9'h0AE;
w_real[635] = 9'h146; w_imag[635] = 9'h0AF;
w_real[636] = 9'h147; w_imag[636] = 9'h0B0;
w_real[637] = 9'h148; w_imag[637] = 9'h0B1;
w_real[638] = 9'h149; w_imag[638] = 9'h0B2;
w_real[639] = 9'h14A; w_imag[639] = 9'h0B3;
w_real[640] = 9'h14B; w_imag[640] = 9'h0B5;
w_real[641] = 9'h14D; w_imag[641] = 9'h0B6;
w_real[642] = 9'h14E; w_imag[642] = 9'h0B7;
w_real[643] = 9'h14F; w_imag[643] = 9'h0B8;
w_real[644] = 9'h150; w_imag[644] = 9'h0B9;
w_real[645] = 9'h151; w_imag[645] = 9'h0BA;
w_real[646] = 9'h152; w_imag[646] = 9'h0BB;
w_real[647] = 9'h153; w_imag[647] = 9'h0BC;
w_real[648] = 9'h155; w_imag[648] = 9'h0BD;
w_real[649] = 9'h156; w_imag[649] = 9'h0BE;
w_real[650] = 9'h157; w_imag[650] = 9'h0BF;
w_real[651] = 9'h158; w_imag[651] = 9'h0C0;
w_real[652] = 9'h159; w_imag[652] = 9'h0C1;
w_real[653] = 9'h15A; w_imag[653] = 9'h0C2;
w_real[654] = 9'h15C; w_imag[654] = 9'h0C3;
w_real[655] = 9'h15D; w_imag[655] = 9'h0C4;
w_real[656] = 9'h15E; w_imag[656] = 9'h0C5;
w_real[657] = 9'h15F; w_imag[657] = 9'h0C6;
w_real[658] = 9'h161; w_imag[658] = 9'h0C7;
w_real[659] = 9'h162; w_imag[659] = 9'h0C8;
w_real[660] = 9'h163; w_imag[660] = 9'h0C9;
w_real[661] = 9'h164; w_imag[661] = 9'h0CA;
w_real[662] = 9'h165; w_imag[662] = 9'h0CB;
w_real[663] = 9'h167; w_imag[663] = 9'h0CC;
w_real[664] = 9'h168; w_imag[664] = 9'h0CD;
w_real[665] = 9'h169; w_imag[665] = 9'h0CE;
w_real[666] = 9'h16B; w_imag[666] = 9'h0CF;
w_real[667] = 9'h16C; w_imag[667] = 9'h0D0;
w_real[668] = 9'h16D; w_imag[668] = 9'h0D1;
w_real[669] = 9'h16E; w_imag[669] = 9'h0D2;
w_real[670] = 9'h170; w_imag[670] = 9'h0D3;
w_real[671] = 9'h171; w_imag[671] = 9'h0D3;
w_real[672] = 9'h172; w_imag[672] = 9'h0D4;
w_real[673] = 9'h174; w_imag[673] = 9'h0D5;
w_real[674] = 9'h175; w_imag[674] = 9'h0D6;
w_real[675] = 9'h176; w_imag[675] = 9'h0D7;
w_real[676] = 9'h178; w_imag[676] = 9'h0D8;
w_real[677] = 9'h179; w_imag[677] = 9'h0D9;
w_real[678] = 9'h17A; w_imag[678] = 9'h0D9;
w_real[679] = 9'h17C; w_imag[679] = 9'h0DA;
w_real[680] = 9'h17D; w_imag[680] = 9'h0DB;
w_real[681] = 9'h17E; w_imag[681] = 9'h0DC;
w_real[682] = 9'h180; w_imag[682] = 9'h0DD;
w_real[683] = 9'h181; w_imag[683] = 9'h0DD;
w_real[684] = 9'h182; w_imag[684] = 9'h0DE;
w_real[685] = 9'h184; w_imag[685] = 9'h0DF;
w_real[686] = 9'h185; w_imag[686] = 9'h0E0;
w_real[687] = 9'h186; w_imag[687] = 9'h0E1;
w_real[688] = 9'h188; w_imag[688] = 9'h0E1;
w_real[689] = 9'h189; w_imag[689] = 9'h0E2;
w_real[690] = 9'h18B; w_imag[690] = 9'h0E3;
w_real[691] = 9'h18C; w_imag[691] = 9'h0E3;
w_real[692] = 9'h18D; w_imag[692] = 9'h0E4;
w_real[693] = 9'h18F; w_imag[693] = 9'h0E5;
w_real[694] = 9'h190; w_imag[694] = 9'h0E6;
w_real[695] = 9'h192; w_imag[695] = 9'h0E6;
w_real[696] = 9'h193; w_imag[696] = 9'h0E7;
w_real[697] = 9'h194; w_imag[697] = 9'h0E8;
w_real[698] = 9'h196; w_imag[698] = 9'h0E8;
w_real[699] = 9'h197; w_imag[699] = 9'h0E9;
w_real[700] = 9'h199; w_imag[700] = 9'h0EA;
w_real[701] = 9'h19A; w_imag[701] = 9'h0EA;
w_real[702] = 9'h19C; w_imag[702] = 9'h0EB;
w_real[703] = 9'h19D; w_imag[703] = 9'h0EB;
w_real[704] = 9'h19F; w_imag[704] = 9'h0EC;
w_real[705] = 9'h1A0; w_imag[705] = 9'h0ED;
w_real[706] = 9'h1A1; w_imag[706] = 9'h0ED;
w_real[707] = 9'h1A3; w_imag[707] = 9'h0EE;
w_real[708] = 9'h1A4; w_imag[708] = 9'h0EE;
w_real[709] = 9'h1A6; w_imag[709] = 9'h0EF;
w_real[710] = 9'h1A7; w_imag[710] = 9'h0EF;
w_real[711] = 9'h1A9; w_imag[711] = 9'h0F0;
w_real[712] = 9'h1AA; w_imag[712] = 9'h0F1;
w_real[713] = 9'h1AC; w_imag[713] = 9'h0F1;
w_real[714] = 9'h1AD; w_imag[714] = 9'h0F2;
w_real[715] = 9'h1AF; w_imag[715] = 9'h0F2;
w_real[716] = 9'h1B0; w_imag[716] = 9'h0F3;
w_real[717] = 9'h1B2; w_imag[717] = 9'h0F3;
w_real[718] = 9'h1B3; w_imag[718] = 9'h0F4;
w_real[719] = 9'h1B5; w_imag[719] = 9'h0F4;
w_real[720] = 9'h1B6; w_imag[720] = 9'h0F4;
w_real[721] = 9'h1B8; w_imag[721] = 9'h0F5;
w_real[722] = 9'h1B9; w_imag[722] = 9'h0F5;
w_real[723] = 9'h1BB; w_imag[723] = 9'h0F6;
w_real[724] = 9'h1BC; w_imag[724] = 9'h0F6;
w_real[725] = 9'h1BE; w_imag[725] = 9'h0F7;
w_real[726] = 9'h1BF; w_imag[726] = 9'h0F7;
w_real[727] = 9'h1C1; w_imag[727] = 9'h0F7;
w_real[728] = 9'h1C2; w_imag[728] = 9'h0F8;
w_real[729] = 9'h1C4; w_imag[729] = 9'h0F8;
w_real[730] = 9'h1C5; w_imag[730] = 9'h0F9;
w_real[731] = 9'h1C7; w_imag[731] = 9'h0F9;
w_real[732] = 9'h1C8; w_imag[732] = 9'h0F9;
w_real[733] = 9'h1CA; w_imag[733] = 9'h0FA;
w_real[734] = 9'h1CB; w_imag[734] = 9'h0FA;
w_real[735] = 9'h1CD; w_imag[735] = 9'h0FA;
w_real[736] = 9'h1CF; w_imag[736] = 9'h0FB;
w_real[737] = 9'h1D0; w_imag[737] = 9'h0FB;
w_real[738] = 9'h1D2; w_imag[738] = 9'h0FB;
w_real[739] = 9'h1D3; w_imag[739] = 9'h0FB;
w_real[740] = 9'h1D5; w_imag[740] = 9'h0FC;
w_real[741] = 9'h1D6; w_imag[741] = 9'h0FC;
w_real[742] = 9'h1D8; w_imag[742] = 9'h0FC;
w_real[743] = 9'h1D9; w_imag[743] = 9'h0FC;
w_real[744] = 9'h1DB; w_imag[744] = 9'h0FD;
w_real[745] = 9'h1DC; w_imag[745] = 9'h0FD;
w_real[746] = 9'h1DE; w_imag[746] = 9'h0FD;
w_real[747] = 9'h1E0; w_imag[747] = 9'h0FD;
w_real[748] = 9'h1E1; w_imag[748] = 9'h0FE;
w_real[749] = 9'h1E3; w_imag[749] = 9'h0FE;
w_real[750] = 9'h1E4; w_imag[750] = 9'h0FE;
w_real[751] = 9'h1E6; w_imag[751] = 9'h0FE;
w_real[752] = 9'h1E7; w_imag[752] = 9'h0FE;
w_real[753] = 9'h1E9; w_imag[753] = 9'h0FE;
w_real[754] = 9'h1EB; w_imag[754] = 9'h0FF;
w_real[755] = 9'h1EC; w_imag[755] = 9'h0FF;
w_real[756] = 9'h1EE; w_imag[756] = 9'h0FF;
w_real[757] = 9'h1EF; w_imag[757] = 9'h0FF;
w_real[758] = 9'h1F1; w_imag[758] = 9'h0FF;
w_real[759] = 9'h1F2; w_imag[759] = 9'h0FF;
w_real[760] = 9'h1F4; w_imag[760] = 9'h0FF;
w_real[761] = 9'h1F6; w_imag[761] = 9'h0FF;
w_real[762] = 9'h1F7; w_imag[762] = 9'h0FF;
w_real[763] = 9'h1F9; w_imag[763] = 9'h0FF;
w_real[764] = 9'h1FA; w_imag[764] = 9'h0FF;
w_real[765] = 9'h1FC; w_imag[765] = 9'h0FF;
w_real[766] = 9'h1FD; w_imag[766] = 9'h0FF;
w_real[767] = 9'h1FF; w_imag[767] = 9'h0FF;
w_real[768] = 9'h000; w_imag[768] = 9'h0FF;
w_real[769] = 9'h001; w_imag[769] = 9'h0FF;
w_real[770] = 9'h003; w_imag[770] = 9'h0FF;
w_real[771] = 9'h004; w_imag[771] = 9'h0FF;
w_real[772] = 9'h006; w_imag[772] = 9'h0FF;
w_real[773] = 9'h007; w_imag[773] = 9'h0FF;
w_real[774] = 9'h009; w_imag[774] = 9'h0FF;
w_real[775] = 9'h00A; w_imag[775] = 9'h0FF;
w_real[776] = 9'h00C; w_imag[776] = 9'h0FF;
w_real[777] = 9'h00E; w_imag[777] = 9'h0FF;
w_real[778] = 9'h00F; w_imag[778] = 9'h0FF;
w_real[779] = 9'h011; w_imag[779] = 9'h0FF;
w_real[780] = 9'h012; w_imag[780] = 9'h0FF;
w_real[781] = 9'h014; w_imag[781] = 9'h0FF;
w_real[782] = 9'h015; w_imag[782] = 9'h0FF;
w_real[783] = 9'h017; w_imag[783] = 9'h0FE;
w_real[784] = 9'h019; w_imag[784] = 9'h0FE;
w_real[785] = 9'h01A; w_imag[785] = 9'h0FE;
w_real[786] = 9'h01C; w_imag[786] = 9'h0FE;
w_real[787] = 9'h01D; w_imag[787] = 9'h0FE;
w_real[788] = 9'h01F; w_imag[788] = 9'h0FE;
w_real[789] = 9'h020; w_imag[789] = 9'h0FD;
w_real[790] = 9'h022; w_imag[790] = 9'h0FD;
w_real[791] = 9'h024; w_imag[791] = 9'h0FD;
w_real[792] = 9'h025; w_imag[792] = 9'h0FD;
w_real[793] = 9'h027; w_imag[793] = 9'h0FC;
w_real[794] = 9'h028; w_imag[794] = 9'h0FC;
w_real[795] = 9'h02A; w_imag[795] = 9'h0FC;
w_real[796] = 9'h02B; w_imag[796] = 9'h0FC;
w_real[797] = 9'h02D; w_imag[797] = 9'h0FB;
w_real[798] = 9'h02E; w_imag[798] = 9'h0FB;
w_real[799] = 9'h030; w_imag[799] = 9'h0FB;
w_real[800] = 9'h031; w_imag[800] = 9'h0FB;
w_real[801] = 9'h033; w_imag[801] = 9'h0FA;
w_real[802] = 9'h035; w_imag[802] = 9'h0FA;
w_real[803] = 9'h036; w_imag[803] = 9'h0FA;
w_real[804] = 9'h038; w_imag[804] = 9'h0F9;
w_real[805] = 9'h039; w_imag[805] = 9'h0F9;
w_real[806] = 9'h03B; w_imag[806] = 9'h0F9;
w_real[807] = 9'h03C; w_imag[807] = 9'h0F8;
w_real[808] = 9'h03E; w_imag[808] = 9'h0F8;
w_real[809] = 9'h03F; w_imag[809] = 9'h0F7;
w_real[810] = 9'h041; w_imag[810] = 9'h0F7;
w_real[811] = 9'h042; w_imag[811] = 9'h0F7;
w_real[812] = 9'h044; w_imag[812] = 9'h0F6;
w_real[813] = 9'h045; w_imag[813] = 9'h0F6;
w_real[814] = 9'h047; w_imag[814] = 9'h0F5;
w_real[815] = 9'h048; w_imag[815] = 9'h0F5;
w_real[816] = 9'h04A; w_imag[816] = 9'h0F4;
w_real[817] = 9'h04B; w_imag[817] = 9'h0F4;
w_real[818] = 9'h04D; w_imag[818] = 9'h0F4;
w_real[819] = 9'h04E; w_imag[819] = 9'h0F3;
w_real[820] = 9'h050; w_imag[820] = 9'h0F3;
w_real[821] = 9'h051; w_imag[821] = 9'h0F2;
w_real[822] = 9'h053; w_imag[822] = 9'h0F2;
w_real[823] = 9'h054; w_imag[823] = 9'h0F1;
w_real[824] = 9'h056; w_imag[824] = 9'h0F1;
w_real[825] = 9'h057; w_imag[825] = 9'h0F0;
w_real[826] = 9'h059; w_imag[826] = 9'h0EF;
w_real[827] = 9'h05A; w_imag[827] = 9'h0EF;
w_real[828] = 9'h05C; w_imag[828] = 9'h0EE;
w_real[829] = 9'h05D; w_imag[829] = 9'h0EE;
w_real[830] = 9'h05F; w_imag[830] = 9'h0ED;
w_real[831] = 9'h060; w_imag[831] = 9'h0ED;
w_real[832] = 9'h061; w_imag[832] = 9'h0EC;
w_real[833] = 9'h063; w_imag[833] = 9'h0EB;
w_real[834] = 9'h064; w_imag[834] = 9'h0EB;
w_real[835] = 9'h066; w_imag[835] = 9'h0EA;
w_real[836] = 9'h067; w_imag[836] = 9'h0EA;
w_real[837] = 9'h069; w_imag[837] = 9'h0E9;
w_real[838] = 9'h06A; w_imag[838] = 9'h0E8;
w_real[839] = 9'h06C; w_imag[839] = 9'h0E8;
w_real[840] = 9'h06D; w_imag[840] = 9'h0E7;
w_real[841] = 9'h06E; w_imag[841] = 9'h0E6;
w_real[842] = 9'h070; w_imag[842] = 9'h0E6;
w_real[843] = 9'h071; w_imag[843] = 9'h0E5;
w_real[844] = 9'h073; w_imag[844] = 9'h0E4;
w_real[845] = 9'h074; w_imag[845] = 9'h0E3;
w_real[846] = 9'h075; w_imag[846] = 9'h0E3;
w_real[847] = 9'h077; w_imag[847] = 9'h0E2;
w_real[848] = 9'h078; w_imag[848] = 9'h0E1;
w_real[849] = 9'h07A; w_imag[849] = 9'h0E1;
w_real[850] = 9'h07B; w_imag[850] = 9'h0E0;
w_real[851] = 9'h07C; w_imag[851] = 9'h0DF;
w_real[852] = 9'h07E; w_imag[852] = 9'h0DE;
w_real[853] = 9'h07F; w_imag[853] = 9'h0DD;
w_real[854] = 9'h080; w_imag[854] = 9'h0DD;
w_real[855] = 9'h082; w_imag[855] = 9'h0DC;
w_real[856] = 9'h083; w_imag[856] = 9'h0DB;
w_real[857] = 9'h084; w_imag[857] = 9'h0DA;
w_real[858] = 9'h086; w_imag[858] = 9'h0D9;
w_real[859] = 9'h087; w_imag[859] = 9'h0D9;
w_real[860] = 9'h088; w_imag[860] = 9'h0D8;
w_real[861] = 9'h08A; w_imag[861] = 9'h0D7;
w_real[862] = 9'h08B; w_imag[862] = 9'h0D6;
w_real[863] = 9'h08C; w_imag[863] = 9'h0D5;
w_real[864] = 9'h08E; w_imag[864] = 9'h0D4;
w_real[865] = 9'h08F; w_imag[865] = 9'h0D3;
w_real[866] = 9'h090; w_imag[866] = 9'h0D3;
w_real[867] = 9'h092; w_imag[867] = 9'h0D2;
w_real[868] = 9'h093; w_imag[868] = 9'h0D1;
w_real[869] = 9'h094; w_imag[869] = 9'h0D0;
w_real[870] = 9'h095; w_imag[870] = 9'h0CF;
w_real[871] = 9'h097; w_imag[871] = 9'h0CE;
w_real[872] = 9'h098; w_imag[872] = 9'h0CD;
w_real[873] = 9'h099; w_imag[873] = 9'h0CC;
w_real[874] = 9'h09B; w_imag[874] = 9'h0CB;
w_real[875] = 9'h09C; w_imag[875] = 9'h0CA;
w_real[876] = 9'h09D; w_imag[876] = 9'h0C9;
w_real[877] = 9'h09E; w_imag[877] = 9'h0C8;
w_real[878] = 9'h09F; w_imag[878] = 9'h0C7;
w_real[879] = 9'h0A1; w_imag[879] = 9'h0C6;
w_real[880] = 9'h0A2; w_imag[880] = 9'h0C5;
w_real[881] = 9'h0A3; w_imag[881] = 9'h0C4;
w_real[882] = 9'h0A4; w_imag[882] = 9'h0C3;
w_real[883] = 9'h0A6; w_imag[883] = 9'h0C2;
w_real[884] = 9'h0A7; w_imag[884] = 9'h0C1;
w_real[885] = 9'h0A8; w_imag[885] = 9'h0C0;
w_real[886] = 9'h0A9; w_imag[886] = 9'h0BF;
w_real[887] = 9'h0AA; w_imag[887] = 9'h0BE;
w_real[888] = 9'h0AB; w_imag[888] = 9'h0BD;
w_real[889] = 9'h0AD; w_imag[889] = 9'h0BC;
w_real[890] = 9'h0AE; w_imag[890] = 9'h0BB;
w_real[891] = 9'h0AF; w_imag[891] = 9'h0BA;
w_real[892] = 9'h0B0; w_imag[892] = 9'h0B9;
w_real[893] = 9'h0B1; w_imag[893] = 9'h0B8;
w_real[894] = 9'h0B2; w_imag[894] = 9'h0B7;
w_real[895] = 9'h0B3; w_imag[895] = 9'h0B6;
w_real[896] = 9'h0B5; w_imag[896] = 9'h0B5;
w_real[897] = 9'h0B6; w_imag[897] = 9'h0B3;
w_real[898] = 9'h0B7; w_imag[898] = 9'h0B2;
w_real[899] = 9'h0B8; w_imag[899] = 9'h0B1;
w_real[900] = 9'h0B9; w_imag[900] = 9'h0B0;
w_real[901] = 9'h0BA; w_imag[901] = 9'h0AF;
w_real[902] = 9'h0BB; w_imag[902] = 9'h0AE;
w_real[903] = 9'h0BC; w_imag[903] = 9'h0AD;
w_real[904] = 9'h0BD; w_imag[904] = 9'h0AB;
w_real[905] = 9'h0BE; w_imag[905] = 9'h0AA;
w_real[906] = 9'h0BF; w_imag[906] = 9'h0A9;
w_real[907] = 9'h0C0; w_imag[907] = 9'h0A8;
w_real[908] = 9'h0C1; w_imag[908] = 9'h0A7;
w_real[909] = 9'h0C2; w_imag[909] = 9'h0A6;
w_real[910] = 9'h0C3; w_imag[910] = 9'h0A4;
w_real[911] = 9'h0C4; w_imag[911] = 9'h0A3;
w_real[912] = 9'h0C5; w_imag[912] = 9'h0A2;
w_real[913] = 9'h0C6; w_imag[913] = 9'h0A1;
w_real[914] = 9'h0C7; w_imag[914] = 9'h09F;
w_real[915] = 9'h0C8; w_imag[915] = 9'h09E;
w_real[916] = 9'h0C9; w_imag[916] = 9'h09D;
w_real[917] = 9'h0CA; w_imag[917] = 9'h09C;
w_real[918] = 9'h0CB; w_imag[918] = 9'h09B;
w_real[919] = 9'h0CC; w_imag[919] = 9'h099;
w_real[920] = 9'h0CD; w_imag[920] = 9'h098;
w_real[921] = 9'h0CE; w_imag[921] = 9'h097;
w_real[922] = 9'h0CF; w_imag[922] = 9'h095;
w_real[923] = 9'h0D0; w_imag[923] = 9'h094;
w_real[924] = 9'h0D1; w_imag[924] = 9'h093;
w_real[925] = 9'h0D2; w_imag[925] = 9'h092;
w_real[926] = 9'h0D3; w_imag[926] = 9'h090;
w_real[927] = 9'h0D3; w_imag[927] = 9'h08F;
w_real[928] = 9'h0D4; w_imag[928] = 9'h08E;
w_real[929] = 9'h0D5; w_imag[929] = 9'h08C;
w_real[930] = 9'h0D6; w_imag[930] = 9'h08B;
w_real[931] = 9'h0D7; w_imag[931] = 9'h08A;
w_real[932] = 9'h0D8; w_imag[932] = 9'h088;
w_real[933] = 9'h0D9; w_imag[933] = 9'h087;
w_real[934] = 9'h0D9; w_imag[934] = 9'h086;
w_real[935] = 9'h0DA; w_imag[935] = 9'h084;
w_real[936] = 9'h0DB; w_imag[936] = 9'h083;
w_real[937] = 9'h0DC; w_imag[937] = 9'h082;
w_real[938] = 9'h0DD; w_imag[938] = 9'h080;
w_real[939] = 9'h0DD; w_imag[939] = 9'h07F;
w_real[940] = 9'h0DE; w_imag[940] = 9'h07E;
w_real[941] = 9'h0DF; w_imag[941] = 9'h07C;
w_real[942] = 9'h0E0; w_imag[942] = 9'h07B;
w_real[943] = 9'h0E1; w_imag[943] = 9'h07A;
w_real[944] = 9'h0E1; w_imag[944] = 9'h078;
w_real[945] = 9'h0E2; w_imag[945] = 9'h077;
w_real[946] = 9'h0E3; w_imag[946] = 9'h075;
w_real[947] = 9'h0E3; w_imag[947] = 9'h074;
w_real[948] = 9'h0E4; w_imag[948] = 9'h073;
w_real[949] = 9'h0E5; w_imag[949] = 9'h071;
w_real[950] = 9'h0E6; w_imag[950] = 9'h070;
w_real[951] = 9'h0E6; w_imag[951] = 9'h06E;
w_real[952] = 9'h0E7; w_imag[952] = 9'h06D;
w_real[953] = 9'h0E8; w_imag[953] = 9'h06C;
w_real[954] = 9'h0E8; w_imag[954] = 9'h06A;
w_real[955] = 9'h0E9; w_imag[955] = 9'h069;
w_real[956] = 9'h0EA; w_imag[956] = 9'h067;
w_real[957] = 9'h0EA; w_imag[957] = 9'h066;
w_real[958] = 9'h0EB; w_imag[958] = 9'h064;
w_real[959] = 9'h0EB; w_imag[959] = 9'h063;
w_real[960] = 9'h0EC; w_imag[960] = 9'h061;
w_real[961] = 9'h0ED; w_imag[961] = 9'h060;
w_real[962] = 9'h0ED; w_imag[962] = 9'h05F;
w_real[963] = 9'h0EE; w_imag[963] = 9'h05D;
w_real[964] = 9'h0EE; w_imag[964] = 9'h05C;
w_real[965] = 9'h0EF; w_imag[965] = 9'h05A;
w_real[966] = 9'h0EF; w_imag[966] = 9'h059;
w_real[967] = 9'h0F0; w_imag[967] = 9'h057;
w_real[968] = 9'h0F1; w_imag[968] = 9'h056;
w_real[969] = 9'h0F1; w_imag[969] = 9'h054;
w_real[970] = 9'h0F2; w_imag[970] = 9'h053;
w_real[971] = 9'h0F2; w_imag[971] = 9'h051;
w_real[972] = 9'h0F3; w_imag[972] = 9'h050;
w_real[973] = 9'h0F3; w_imag[973] = 9'h04E;
w_real[974] = 9'h0F4; w_imag[974] = 9'h04D;
w_real[975] = 9'h0F4; w_imag[975] = 9'h04B;
w_real[976] = 9'h0F4; w_imag[976] = 9'h04A;
w_real[977] = 9'h0F5; w_imag[977] = 9'h048;
w_real[978] = 9'h0F5; w_imag[978] = 9'h047;
w_real[979] = 9'h0F6; w_imag[979] = 9'h045;
w_real[980] = 9'h0F6; w_imag[980] = 9'h044;
w_real[981] = 9'h0F7; w_imag[981] = 9'h042;
w_real[982] = 9'h0F7; w_imag[982] = 9'h041;
w_real[983] = 9'h0F7; w_imag[983] = 9'h03F;
w_real[984] = 9'h0F8; w_imag[984] = 9'h03E;
w_real[985] = 9'h0F8; w_imag[985] = 9'h03C;
w_real[986] = 9'h0F9; w_imag[986] = 9'h03B;
w_real[987] = 9'h0F9; w_imag[987] = 9'h039;
w_real[988] = 9'h0F9; w_imag[988] = 9'h038;
w_real[989] = 9'h0FA; w_imag[989] = 9'h036;
w_real[990] = 9'h0FA; w_imag[990] = 9'h035;
w_real[991] = 9'h0FA; w_imag[991] = 9'h033;
w_real[992] = 9'h0FB; w_imag[992] = 9'h031;
w_real[993] = 9'h0FB; w_imag[993] = 9'h030;
w_real[994] = 9'h0FB; w_imag[994] = 9'h02E;
w_real[995] = 9'h0FB; w_imag[995] = 9'h02D;
w_real[996] = 9'h0FC; w_imag[996] = 9'h02B;
w_real[997] = 9'h0FC; w_imag[997] = 9'h02A;
w_real[998] = 9'h0FC; w_imag[998] = 9'h028;
w_real[999] = 9'h0FC; w_imag[999] = 9'h027;
w_real[1000] = 9'h0FD; w_imag[1000] = 9'h025;
w_real[1001] = 9'h0FD; w_imag[1001] = 9'h024;
w_real[1002] = 9'h0FD; w_imag[1002] = 9'h022;
w_real[1003] = 9'h0FD; w_imag[1003] = 9'h020;
w_real[1004] = 9'h0FE; w_imag[1004] = 9'h01F;
w_real[1005] = 9'h0FE; w_imag[1005] = 9'h01D;
w_real[1006] = 9'h0FE; w_imag[1006] = 9'h01C;
w_real[1007] = 9'h0FE; w_imag[1007] = 9'h01A;
w_real[1008] = 9'h0FE; w_imag[1008] = 9'h019;
w_real[1009] = 9'h0FE; w_imag[1009] = 9'h017;
w_real[1010] = 9'h0FF; w_imag[1010] = 9'h015;
w_real[1011] = 9'h0FF; w_imag[1011] = 9'h014;
w_real[1012] = 9'h0FF; w_imag[1012] = 9'h012;
w_real[1013] = 9'h0FF; w_imag[1013] = 9'h011;
w_real[1014] = 9'h0FF; w_imag[1014] = 9'h00F;
w_real[1015] = 9'h0FF; w_imag[1015] = 9'h00E;
w_real[1016] = 9'h0FF; w_imag[1016] = 9'h00C;
w_real[1017] = 9'h0FF; w_imag[1017] = 9'h00A;
w_real[1018] = 9'h0FF; w_imag[1018] = 9'h009;
w_real[1019] = 9'h0FF; w_imag[1019] = 9'h007;
w_real[1020] = 9'h0FF; w_imag[1020] = 9'h006;
w_real[1021] = 9'h0FF; w_imag[1021] = 9'h004;
w_real[1022] = 9'h0FF; w_imag[1022] = 9'h003;
w_real[1023] = 9'h0FF; w_imag[1023] = 9'h001;
