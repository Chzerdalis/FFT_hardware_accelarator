0 0
1419 -7137
8582 -20721
34856 -52166
110556 -110556
-44543 29763
-49000 20296
-42272 8408
-39196 0
-42272 -8408
-49000 -20296
-44543 -29763
110556 110556
34856 52166
8582 20721
1419 7137
