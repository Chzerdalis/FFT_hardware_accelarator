w_real[0] = 9'h0FF; w_imag[0] = 9'h000;
w_real[1] = 9'h0FF; w_imag[1] = 9'h1FA;
w_real[2] = 9'h0FF; w_imag[2] = 9'h1F4;
w_real[3] = 9'h0FF; w_imag[3] = 9'h1EE;
w_real[4] = 9'h0FE; w_imag[4] = 9'h1E7;
w_real[5] = 9'h0FE; w_imag[5] = 9'h1E1;
w_real[6] = 9'h0FD; w_imag[6] = 9'h1DB;
w_real[7] = 9'h0FC; w_imag[7] = 9'h1D5;
w_real[8] = 9'h0FB; w_imag[8] = 9'h1CF;
w_real[9] = 9'h0F9; w_imag[9] = 9'h1C8;
w_real[10] = 9'h0F8; w_imag[10] = 9'h1C2;
w_real[11] = 9'h0F6; w_imag[11] = 9'h1BC;
w_real[12] = 9'h0F4; w_imag[12] = 9'h1B6;
w_real[13] = 9'h0F3; w_imag[13] = 9'h1B0;
w_real[14] = 9'h0F1; w_imag[14] = 9'h1AA;
w_real[15] = 9'h0EE; w_imag[15] = 9'h1A4;
w_real[16] = 9'h0EC; w_imag[16] = 9'h19F;
w_real[17] = 9'h0EA; w_imag[17] = 9'h199;
w_real[18] = 9'h0E7; w_imag[18] = 9'h193;
w_real[19] = 9'h0E4; w_imag[19] = 9'h18D;
w_real[20] = 9'h0E1; w_imag[20] = 9'h188;
w_real[21] = 9'h0DE; w_imag[21] = 9'h182;
w_real[22] = 9'h0DB; w_imag[22] = 9'h17D;
w_real[23] = 9'h0D8; w_imag[23] = 9'h178;
w_real[24] = 9'h0D4; w_imag[24] = 9'h172;
w_real[25] = 9'h0D1; w_imag[25] = 9'h16D;
w_real[26] = 9'h0CD; w_imag[26] = 9'h168;
w_real[27] = 9'h0C9; w_imag[27] = 9'h163;
w_real[28] = 9'h0C5; w_imag[28] = 9'h15E;
w_real[29] = 9'h0C1; w_imag[29] = 9'h159;
w_real[30] = 9'h0BD; w_imag[30] = 9'h155;
w_real[31] = 9'h0B9; w_imag[31] = 9'h150;
w_real[32] = 9'h0B5; w_imag[32] = 9'h14B;
w_real[33] = 9'h0B0; w_imag[33] = 9'h147;
w_real[34] = 9'h0AB; w_imag[34] = 9'h143;
w_real[35] = 9'h0A7; w_imag[35] = 9'h13F;
w_real[36] = 9'h0A2; w_imag[36] = 9'h13B;
w_real[37] = 9'h09D; w_imag[37] = 9'h137;
w_real[38] = 9'h098; w_imag[38] = 9'h133;
w_real[39] = 9'h093; w_imag[39] = 9'h12F;
w_real[40] = 9'h08E; w_imag[40] = 9'h12C;
w_real[41] = 9'h088; w_imag[41] = 9'h128;
w_real[42] = 9'h083; w_imag[42] = 9'h125;
w_real[43] = 9'h07E; w_imag[43] = 9'h122;
w_real[44] = 9'h078; w_imag[44] = 9'h11F;
w_real[45] = 9'h073; w_imag[45] = 9'h11C;
w_real[46] = 9'h06D; w_imag[46] = 9'h119;
w_real[47] = 9'h067; w_imag[47] = 9'h116;
w_real[48] = 9'h061; w_imag[48] = 9'h114;
w_real[49] = 9'h05C; w_imag[49] = 9'h112;
w_real[50] = 9'h056; w_imag[50] = 9'h10F;
w_real[51] = 9'h050; w_imag[51] = 9'h10D;
w_real[52] = 9'h04A; w_imag[52] = 9'h10C;
w_real[53] = 9'h044; w_imag[53] = 9'h10A;
w_real[54] = 9'h03E; w_imag[54] = 9'h108;
w_real[55] = 9'h038; w_imag[55] = 9'h107;
w_real[56] = 9'h031; w_imag[56] = 9'h105;
w_real[57] = 9'h02B; w_imag[57] = 9'h104;
w_real[58] = 9'h025; w_imag[58] = 9'h103;
w_real[59] = 9'h01F; w_imag[59] = 9'h102;
w_real[60] = 9'h019; w_imag[60] = 9'h102;
w_real[61] = 9'h012; w_imag[61] = 9'h101;
w_real[62] = 9'h00C; w_imag[62] = 9'h101;
w_real[63] = 9'h006; w_imag[63] = 9'h101;
w_real[64] = 9'h000; w_imag[64] = 9'h100;
w_real[65] = 9'h1FA; w_imag[65] = 9'h101;
w_real[66] = 9'h1F4; w_imag[66] = 9'h101;
w_real[67] = 9'h1EE; w_imag[67] = 9'h101;
w_real[68] = 9'h1E7; w_imag[68] = 9'h102;
w_real[69] = 9'h1E1; w_imag[69] = 9'h102;
w_real[70] = 9'h1DB; w_imag[70] = 9'h103;
w_real[71] = 9'h1D5; w_imag[71] = 9'h104;
w_real[72] = 9'h1CF; w_imag[72] = 9'h105;
w_real[73] = 9'h1C8; w_imag[73] = 9'h107;
w_real[74] = 9'h1C2; w_imag[74] = 9'h108;
w_real[75] = 9'h1BC; w_imag[75] = 9'h10A;
w_real[76] = 9'h1B6; w_imag[76] = 9'h10C;
w_real[77] = 9'h1B0; w_imag[77] = 9'h10D;
w_real[78] = 9'h1AA; w_imag[78] = 9'h10F;
w_real[79] = 9'h1A4; w_imag[79] = 9'h112;
w_real[80] = 9'h19F; w_imag[80] = 9'h114;
w_real[81] = 9'h199; w_imag[81] = 9'h116;
w_real[82] = 9'h193; w_imag[82] = 9'h119;
w_real[83] = 9'h18D; w_imag[83] = 9'h11C;
w_real[84] = 9'h188; w_imag[84] = 9'h11F;
w_real[85] = 9'h182; w_imag[85] = 9'h122;
w_real[86] = 9'h17D; w_imag[86] = 9'h125;
w_real[87] = 9'h178; w_imag[87] = 9'h128;
w_real[88] = 9'h172; w_imag[88] = 9'h12C;
w_real[89] = 9'h16D; w_imag[89] = 9'h12F;
w_real[90] = 9'h168; w_imag[90] = 9'h133;
w_real[91] = 9'h163; w_imag[91] = 9'h137;
w_real[92] = 9'h15E; w_imag[92] = 9'h13B;
w_real[93] = 9'h159; w_imag[93] = 9'h13F;
w_real[94] = 9'h155; w_imag[94] = 9'h143;
w_real[95] = 9'h150; w_imag[95] = 9'h147;
w_real[96] = 9'h14B; w_imag[96] = 9'h14B;
w_real[97] = 9'h147; w_imag[97] = 9'h150;
w_real[98] = 9'h143; w_imag[98] = 9'h155;
w_real[99] = 9'h13F; w_imag[99] = 9'h159;
w_real[100] = 9'h13B; w_imag[100] = 9'h15E;
w_real[101] = 9'h137; w_imag[101] = 9'h163;
w_real[102] = 9'h133; w_imag[102] = 9'h168;
w_real[103] = 9'h12F; w_imag[103] = 9'h16D;
w_real[104] = 9'h12C; w_imag[104] = 9'h172;
w_real[105] = 9'h128; w_imag[105] = 9'h178;
w_real[106] = 9'h125; w_imag[106] = 9'h17D;
w_real[107] = 9'h122; w_imag[107] = 9'h182;
w_real[108] = 9'h11F; w_imag[108] = 9'h188;
w_real[109] = 9'h11C; w_imag[109] = 9'h18D;
w_real[110] = 9'h119; w_imag[110] = 9'h193;
w_real[111] = 9'h116; w_imag[111] = 9'h199;
w_real[112] = 9'h114; w_imag[112] = 9'h19F;
w_real[113] = 9'h112; w_imag[113] = 9'h1A4;
w_real[114] = 9'h10F; w_imag[114] = 9'h1AA;
w_real[115] = 9'h10D; w_imag[115] = 9'h1B0;
w_real[116] = 9'h10C; w_imag[116] = 9'h1B6;
w_real[117] = 9'h10A; w_imag[117] = 9'h1BC;
w_real[118] = 9'h108; w_imag[118] = 9'h1C2;
w_real[119] = 9'h107; w_imag[119] = 9'h1C8;
w_real[120] = 9'h105; w_imag[120] = 9'h1CF;
w_real[121] = 9'h104; w_imag[121] = 9'h1D5;
w_real[122] = 9'h103; w_imag[122] = 9'h1DB;
w_real[123] = 9'h102; w_imag[123] = 9'h1E1;
w_real[124] = 9'h102; w_imag[124] = 9'h1E7;
w_real[125] = 9'h101; w_imag[125] = 9'h1EE;
w_real[126] = 9'h101; w_imag[126] = 9'h1F4;
w_real[127] = 9'h101; w_imag[127] = 9'h1FA;
w_real[128] = 9'h100; w_imag[128] = 9'h000;
w_real[129] = 9'h101; w_imag[129] = 9'h006;
w_real[130] = 9'h101; w_imag[130] = 9'h00C;
w_real[131] = 9'h101; w_imag[131] = 9'h012;
w_real[132] = 9'h102; w_imag[132] = 9'h019;
w_real[133] = 9'h102; w_imag[133] = 9'h01F;
w_real[134] = 9'h103; w_imag[134] = 9'h025;
w_real[135] = 9'h104; w_imag[135] = 9'h02B;
w_real[136] = 9'h105; w_imag[136] = 9'h031;
w_real[137] = 9'h107; w_imag[137] = 9'h038;
w_real[138] = 9'h108; w_imag[138] = 9'h03E;
w_real[139] = 9'h10A; w_imag[139] = 9'h044;
w_real[140] = 9'h10C; w_imag[140] = 9'h04A;
w_real[141] = 9'h10D; w_imag[141] = 9'h050;
w_real[142] = 9'h10F; w_imag[142] = 9'h056;
w_real[143] = 9'h112; w_imag[143] = 9'h05C;
w_real[144] = 9'h114; w_imag[144] = 9'h061;
w_real[145] = 9'h116; w_imag[145] = 9'h067;
w_real[146] = 9'h119; w_imag[146] = 9'h06D;
w_real[147] = 9'h11C; w_imag[147] = 9'h073;
w_real[148] = 9'h11F; w_imag[148] = 9'h078;
w_real[149] = 9'h122; w_imag[149] = 9'h07E;
w_real[150] = 9'h125; w_imag[150] = 9'h083;
w_real[151] = 9'h128; w_imag[151] = 9'h088;
w_real[152] = 9'h12C; w_imag[152] = 9'h08E;
w_real[153] = 9'h12F; w_imag[153] = 9'h093;
w_real[154] = 9'h133; w_imag[154] = 9'h098;
w_real[155] = 9'h137; w_imag[155] = 9'h09D;
w_real[156] = 9'h13B; w_imag[156] = 9'h0A2;
w_real[157] = 9'h13F; w_imag[157] = 9'h0A7;
w_real[158] = 9'h143; w_imag[158] = 9'h0AB;
w_real[159] = 9'h147; w_imag[159] = 9'h0B0;
w_real[160] = 9'h14B; w_imag[160] = 9'h0B5;
w_real[161] = 9'h150; w_imag[161] = 9'h0B9;
w_real[162] = 9'h155; w_imag[162] = 9'h0BD;
w_real[163] = 9'h159; w_imag[163] = 9'h0C1;
w_real[164] = 9'h15E; w_imag[164] = 9'h0C5;
w_real[165] = 9'h163; w_imag[165] = 9'h0C9;
w_real[166] = 9'h168; w_imag[166] = 9'h0CD;
w_real[167] = 9'h16D; w_imag[167] = 9'h0D1;
w_real[168] = 9'h172; w_imag[168] = 9'h0D4;
w_real[169] = 9'h178; w_imag[169] = 9'h0D8;
w_real[170] = 9'h17D; w_imag[170] = 9'h0DB;
w_real[171] = 9'h182; w_imag[171] = 9'h0DE;
w_real[172] = 9'h188; w_imag[172] = 9'h0E1;
w_real[173] = 9'h18D; w_imag[173] = 9'h0E4;
w_real[174] = 9'h193; w_imag[174] = 9'h0E7;
w_real[175] = 9'h199; w_imag[175] = 9'h0EA;
w_real[176] = 9'h19F; w_imag[176] = 9'h0EC;
w_real[177] = 9'h1A4; w_imag[177] = 9'h0EE;
w_real[178] = 9'h1AA; w_imag[178] = 9'h0F1;
w_real[179] = 9'h1B0; w_imag[179] = 9'h0F3;
w_real[180] = 9'h1B6; w_imag[180] = 9'h0F4;
w_real[181] = 9'h1BC; w_imag[181] = 9'h0F6;
w_real[182] = 9'h1C2; w_imag[182] = 9'h0F8;
w_real[183] = 9'h1C8; w_imag[183] = 9'h0F9;
w_real[184] = 9'h1CF; w_imag[184] = 9'h0FB;
w_real[185] = 9'h1D5; w_imag[185] = 9'h0FC;
w_real[186] = 9'h1DB; w_imag[186] = 9'h0FD;
w_real[187] = 9'h1E1; w_imag[187] = 9'h0FE;
w_real[188] = 9'h1E7; w_imag[188] = 9'h0FE;
w_real[189] = 9'h1EE; w_imag[189] = 9'h0FF;
w_real[190] = 9'h1F4; w_imag[190] = 9'h0FF;
w_real[191] = 9'h1FA; w_imag[191] = 9'h0FF;
w_real[192] = 9'h000; w_imag[192] = 9'h0FF;
w_real[193] = 9'h006; w_imag[193] = 9'h0FF;
w_real[194] = 9'h00C; w_imag[194] = 9'h0FF;
w_real[195] = 9'h012; w_imag[195] = 9'h0FF;
w_real[196] = 9'h019; w_imag[196] = 9'h0FE;
w_real[197] = 9'h01F; w_imag[197] = 9'h0FE;
w_real[198] = 9'h025; w_imag[198] = 9'h0FD;
w_real[199] = 9'h02B; w_imag[199] = 9'h0FC;
w_real[200] = 9'h031; w_imag[200] = 9'h0FB;
w_real[201] = 9'h038; w_imag[201] = 9'h0F9;
w_real[202] = 9'h03E; w_imag[202] = 9'h0F8;
w_real[203] = 9'h044; w_imag[203] = 9'h0F6;
w_real[204] = 9'h04A; w_imag[204] = 9'h0F4;
w_real[205] = 9'h050; w_imag[205] = 9'h0F3;
w_real[206] = 9'h056; w_imag[206] = 9'h0F1;
w_real[207] = 9'h05C; w_imag[207] = 9'h0EE;
w_real[208] = 9'h061; w_imag[208] = 9'h0EC;
w_real[209] = 9'h067; w_imag[209] = 9'h0EA;
w_real[210] = 9'h06D; w_imag[210] = 9'h0E7;
w_real[211] = 9'h073; w_imag[211] = 9'h0E4;
w_real[212] = 9'h078; w_imag[212] = 9'h0E1;
w_real[213] = 9'h07E; w_imag[213] = 9'h0DE;
w_real[214] = 9'h083; w_imag[214] = 9'h0DB;
w_real[215] = 9'h088; w_imag[215] = 9'h0D8;
w_real[216] = 9'h08E; w_imag[216] = 9'h0D4;
w_real[217] = 9'h093; w_imag[217] = 9'h0D1;
w_real[218] = 9'h098; w_imag[218] = 9'h0CD;
w_real[219] = 9'h09D; w_imag[219] = 9'h0C9;
w_real[220] = 9'h0A2; w_imag[220] = 9'h0C5;
w_real[221] = 9'h0A7; w_imag[221] = 9'h0C1;
w_real[222] = 9'h0AB; w_imag[222] = 9'h0BD;
w_real[223] = 9'h0B0; w_imag[223] = 9'h0B9;
w_real[224] = 9'h0B5; w_imag[224] = 9'h0B5;
w_real[225] = 9'h0B9; w_imag[225] = 9'h0B0;
w_real[226] = 9'h0BD; w_imag[226] = 9'h0AB;
w_real[227] = 9'h0C1; w_imag[227] = 9'h0A7;
w_real[228] = 9'h0C5; w_imag[228] = 9'h0A2;
w_real[229] = 9'h0C9; w_imag[229] = 9'h09D;
w_real[230] = 9'h0CD; w_imag[230] = 9'h098;
w_real[231] = 9'h0D1; w_imag[231] = 9'h093;
w_real[232] = 9'h0D4; w_imag[232] = 9'h08E;
w_real[233] = 9'h0D8; w_imag[233] = 9'h088;
w_real[234] = 9'h0DB; w_imag[234] = 9'h083;
w_real[235] = 9'h0DE; w_imag[235] = 9'h07E;
w_real[236] = 9'h0E1; w_imag[236] = 9'h078;
w_real[237] = 9'h0E4; w_imag[237] = 9'h073;
w_real[238] = 9'h0E7; w_imag[238] = 9'h06D;
w_real[239] = 9'h0EA; w_imag[239] = 9'h067;
w_real[240] = 9'h0EC; w_imag[240] = 9'h061;
w_real[241] = 9'h0EE; w_imag[241] = 9'h05C;
w_real[242] = 9'h0F1; w_imag[242] = 9'h056;
w_real[243] = 9'h0F3; w_imag[243] = 9'h050;
w_real[244] = 9'h0F4; w_imag[244] = 9'h04A;
w_real[245] = 9'h0F6; w_imag[245] = 9'h044;
w_real[246] = 9'h0F8; w_imag[246] = 9'h03E;
w_real[247] = 9'h0F9; w_imag[247] = 9'h038;
w_real[248] = 9'h0FB; w_imag[248] = 9'h031;
w_real[249] = 9'h0FC; w_imag[249] = 9'h02B;
w_real[250] = 9'h0FD; w_imag[250] = 9'h025;
w_real[251] = 9'h0FE; w_imag[251] = 9'h01F;
w_real[252] = 9'h0FE; w_imag[252] = 9'h019;
w_real[253] = 9'h0FF; w_imag[253] = 9'h012;
w_real[254] = 9'h0FF; w_imag[254] = 9'h00C;
w_real[255] = 9'h0FF; w_imag[255] = 9'h006;
