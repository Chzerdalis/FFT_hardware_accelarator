w_real[0] = 16'h7FFF; w_imag[0] = 16'h0000;
w_real[1] = 16'h7FFF; w_imag[1] = 16'hFF37;
w_real[2] = 16'h7FFD; w_imag[2] = 16'hFE6E;
w_real[3] = 16'h7FFA; w_imag[3] = 16'hFDA5;
w_real[4] = 16'h7FF6; w_imag[4] = 16'hFCDC;
w_real[5] = 16'h7FF0; w_imag[5] = 16'hFC13;
w_real[6] = 16'h7FE9; w_imag[6] = 16'hFB4A;
w_real[7] = 16'h7FE1; w_imag[7] = 16'hFA81;
w_real[8] = 16'h7FD8; w_imag[8] = 16'hF9B9;
w_real[9] = 16'h7FCE; w_imag[9] = 16'hF8F0;
w_real[10] = 16'h7FC2; w_imag[10] = 16'hF827;
w_real[11] = 16'h7FB5; w_imag[11] = 16'hF75E;
w_real[12] = 16'h7FA7; w_imag[12] = 16'hF696;
w_real[13] = 16'h7F97; w_imag[13] = 16'hF5CD;
w_real[14] = 16'h7F87; w_imag[14] = 16'hF505;
w_real[15] = 16'h7F75; w_imag[15] = 16'hF43D;
w_real[16] = 16'h7F62; w_imag[16] = 16'hF375;
w_real[17] = 16'h7F4D; w_imag[17] = 16'hF2AD;
w_real[18] = 16'h7F38; w_imag[18] = 16'hF1E5;
w_real[19] = 16'h7F21; w_imag[19] = 16'hF11D;
w_real[20] = 16'h7F09; w_imag[20] = 16'hF055;
w_real[21] = 16'h7EF0; w_imag[21] = 16'hEF8E;
w_real[22] = 16'h7ED5; w_imag[22] = 16'hEEC7;
w_real[23] = 16'h7EBA; w_imag[23] = 16'hEDFF;
w_real[24] = 16'h7E9D; w_imag[24] = 16'hED38;
w_real[25] = 16'h7E7F; w_imag[25] = 16'hEC72;
w_real[26] = 16'h7E5F; w_imag[26] = 16'hEBAB;
w_real[27] = 16'h7E3F; w_imag[27] = 16'hEAE5;
w_real[28] = 16'h7E1D; w_imag[28] = 16'hEA1E;
w_real[29] = 16'h7DFA; w_imag[29] = 16'hE958;
w_real[30] = 16'h7DD6; w_imag[30] = 16'hE893;
w_real[31] = 16'h7DB0; w_imag[31] = 16'hE7CD;
w_real[32] = 16'h7D8A; w_imag[32] = 16'hE708;
w_real[33] = 16'h7D62; w_imag[33] = 16'hE643;
w_real[34] = 16'h7D39; w_imag[34] = 16'hE57E;
w_real[35] = 16'h7D0F; w_imag[35] = 16'hE4B9;
w_real[36] = 16'h7CE3; w_imag[36] = 16'hE3F5;
w_real[37] = 16'h7CB7; w_imag[37] = 16'hE331;
w_real[38] = 16'h7C89; w_imag[38] = 16'hE26D;
w_real[39] = 16'h7C5A; w_imag[39] = 16'hE1AA;
w_real[40] = 16'h7C29; w_imag[40] = 16'hE0E7;
w_real[41] = 16'h7BF8; w_imag[41] = 16'hE024;
w_real[42] = 16'h7BC5; w_imag[42] = 16'hDF61;
w_real[43] = 16'h7B92; w_imag[43] = 16'hDE9F;
w_real[44] = 16'h7B5D; w_imag[44] = 16'hDDDD;
w_real[45] = 16'h7B26; w_imag[45] = 16'hDD1B;
w_real[46] = 16'h7AEF; w_imag[46] = 16'hDC5A;
w_real[47] = 16'h7AB6; w_imag[47] = 16'hDB99;
w_real[48] = 16'h7A7D; w_imag[48] = 16'hDAD8;
w_real[49] = 16'h7A42; w_imag[49] = 16'hDA18;
w_real[50] = 16'h7A05; w_imag[50] = 16'hD958;
w_real[51] = 16'h79C8; w_imag[51] = 16'hD899;
w_real[52] = 16'h798A; w_imag[52] = 16'hD7DA;
w_real[53] = 16'h794A; w_imag[53] = 16'hD71B;
w_real[54] = 16'h7909; w_imag[54] = 16'hD65D;
w_real[55] = 16'h78C7; w_imag[55] = 16'hD59F;
w_real[56] = 16'h7884; w_imag[56] = 16'hD4E1;
w_real[57] = 16'h7840; w_imag[57] = 16'hD424;
w_real[58] = 16'h77FA; w_imag[58] = 16'hD368;
w_real[59] = 16'h77B4; w_imag[59] = 16'hD2AB;
w_real[60] = 16'h776C; w_imag[60] = 16'hD1EF;
w_real[61] = 16'h7723; w_imag[61] = 16'hD134;
w_real[62] = 16'h76D9; w_imag[62] = 16'hD079;
w_real[63] = 16'h768E; w_imag[63] = 16'hCFBF;
w_real[64] = 16'h7641; w_imag[64] = 16'hCF05;
w_real[65] = 16'h75F4; w_imag[65] = 16'hCE4B;
w_real[66] = 16'h75A5; w_imag[66] = 16'hCD92;
w_real[67] = 16'h7555; w_imag[67] = 16'hCCDA;
w_real[68] = 16'h7504; w_imag[68] = 16'hCC22;
w_real[69] = 16'h74B2; w_imag[69] = 16'hCB6A;
w_real[70] = 16'h745F; w_imag[70] = 16'hCAB3;
w_real[71] = 16'h740B; w_imag[71] = 16'hC9FC;
w_real[72] = 16'h73B5; w_imag[72] = 16'hC946;
w_real[73] = 16'h735F; w_imag[73] = 16'hC891;
w_real[74] = 16'h7307; w_imag[74] = 16'hC7DC;
w_real[75] = 16'h72AF; w_imag[75] = 16'hC728;
w_real[76] = 16'h7255; w_imag[76] = 16'hC674;
w_real[77] = 16'h71FA; w_imag[77] = 16'hC5C0;
w_real[78] = 16'h719E; w_imag[78] = 16'hC50E;
w_real[79] = 16'h7141; w_imag[79] = 16'hC45B;
w_real[80] = 16'h70E2; w_imag[80] = 16'hC3AA;
w_real[81] = 16'h7083; w_imag[81] = 16'hC2F9;
w_real[82] = 16'h7023; w_imag[82] = 16'hC248;
w_real[83] = 16'h6FC1; w_imag[83] = 16'hC198;
w_real[84] = 16'h6F5F; w_imag[84] = 16'hC0E9;
w_real[85] = 16'h6EFB; w_imag[85] = 16'hC03B;
w_real[86] = 16'h6E96; w_imag[86] = 16'hBF8D;
w_real[87] = 16'h6E30; w_imag[87] = 16'hBEDF;
w_real[88] = 16'h6DCA; w_imag[88] = 16'hBE32;
w_real[89] = 16'h6D62; w_imag[89] = 16'hBD86;
w_real[90] = 16'h6CF9; w_imag[90] = 16'hBCDB;
w_real[91] = 16'h6C8F; w_imag[91] = 16'hBC30;
w_real[92] = 16'h6C24; w_imag[92] = 16'hBB86;
w_real[93] = 16'h6BB8; w_imag[93] = 16'hBADC;
w_real[94] = 16'h6B4A; w_imag[94] = 16'hBA33;
w_real[95] = 16'h6ADC; w_imag[95] = 16'hB98B;
w_real[96] = 16'h6A6D; w_imag[96] = 16'hB8E4;
w_real[97] = 16'h69FD; w_imag[97] = 16'hB83D;
w_real[98] = 16'h698C; w_imag[98] = 16'hB797;
w_real[99] = 16'h6919; w_imag[99] = 16'hB6F1;
w_real[100] = 16'h68A6; w_imag[100] = 16'hB64C;
w_real[101] = 16'h6832; w_imag[101] = 16'hB5A8;
w_real[102] = 16'h67BD; w_imag[102] = 16'hB505;
w_real[103] = 16'h6746; w_imag[103] = 16'hB462;
w_real[104] = 16'h66CF; w_imag[104] = 16'hB3C1;
w_real[105] = 16'h6657; w_imag[105] = 16'hB31F;
w_real[106] = 16'h65DD; w_imag[106] = 16'hB27F;
w_real[107] = 16'h6563; w_imag[107] = 16'hB1DF;
w_real[108] = 16'h64E8; w_imag[108] = 16'hB141;
w_real[109] = 16'h646C; w_imag[109] = 16'hB0A2;
w_real[110] = 16'h63EF; w_imag[110] = 16'hB005;
w_real[111] = 16'h6371; w_imag[111] = 16'hAF69;
w_real[112] = 16'h62F2; w_imag[112] = 16'hAECD;
w_real[113] = 16'h6271; w_imag[113] = 16'hAE32;
w_real[114] = 16'h61F1; w_imag[114] = 16'hAD97;
w_real[115] = 16'h616F; w_imag[115] = 16'hACFE;
w_real[116] = 16'h60EC; w_imag[116] = 16'hAC65;
w_real[117] = 16'h6068; w_imag[117] = 16'hABCD;
w_real[118] = 16'h5FE3; w_imag[118] = 16'hAB36;
w_real[119] = 16'h5F5E; w_imag[119] = 16'hAAA0;
w_real[120] = 16'h5ED7; w_imag[120] = 16'hAA0B;
w_real[121] = 16'h5E50; w_imag[121] = 16'hA976;
w_real[122] = 16'h5DC7; w_imag[122] = 16'hA8E3;
w_real[123] = 16'h5D3E; w_imag[123] = 16'hA850;
w_real[124] = 16'h5CB4; w_imag[124] = 16'hA7BE;
w_real[125] = 16'h5C29; w_imag[125] = 16'hA72C;
w_real[126] = 16'h5B9D; w_imag[126] = 16'hA69C;
w_real[127] = 16'h5B10; w_imag[127] = 16'hA60D;
w_real[128] = 16'h5A82; w_imag[128] = 16'hA57E;
w_real[129] = 16'h59F3; w_imag[129] = 16'hA4F0;
w_real[130] = 16'h5964; w_imag[130] = 16'hA463;
w_real[131] = 16'h58D4; w_imag[131] = 16'hA3D7;
w_real[132] = 16'h5842; w_imag[132] = 16'hA34C;
w_real[133] = 16'h57B0; w_imag[133] = 16'hA2C2;
w_real[134] = 16'h571D; w_imag[134] = 16'hA239;
w_real[135] = 16'h568A; w_imag[135] = 16'hA1B0;
w_real[136] = 16'h55F5; w_imag[136] = 16'hA129;
w_real[137] = 16'h5560; w_imag[137] = 16'hA0A2;
w_real[138] = 16'h54CA; w_imag[138] = 16'hA01D;
w_real[139] = 16'h5433; w_imag[139] = 16'h9F98;
w_real[140] = 16'h539B; w_imag[140] = 16'h9F14;
w_real[141] = 16'h5302; w_imag[141] = 16'h9E91;
w_real[142] = 16'h5269; w_imag[142] = 16'h9E0F;
w_real[143] = 16'h51CE; w_imag[143] = 16'h9D8F;
w_real[144] = 16'h5133; w_imag[144] = 16'h9D0E;
w_real[145] = 16'h5097; w_imag[145] = 16'h9C8F;
w_real[146] = 16'h4FFB; w_imag[146] = 16'h9C11;
w_real[147] = 16'h4F5E; w_imag[147] = 16'h9B94;
w_real[148] = 16'h4EBF; w_imag[148] = 16'h9B18;
w_real[149] = 16'h4E21; w_imag[149] = 16'h9A9D;
w_real[150] = 16'h4D81; w_imag[150] = 16'h9A23;
w_real[151] = 16'h4CE1; w_imag[151] = 16'h99A9;
w_real[152] = 16'h4C3F; w_imag[152] = 16'h9931;
w_real[153] = 16'h4B9E; w_imag[153] = 16'h98BA;
w_real[154] = 16'h4AFB; w_imag[154] = 16'h9843;
w_real[155] = 16'h4A58; w_imag[155] = 16'h97CE;
w_real[156] = 16'h49B4; w_imag[156] = 16'h975A;
w_real[157] = 16'h490F; w_imag[157] = 16'h96E7;
w_real[158] = 16'h4869; w_imag[158] = 16'h9674;
w_real[159] = 16'h47C3; w_imag[159] = 16'h9603;
w_real[160] = 16'h471C; w_imag[160] = 16'h9593;
w_real[161] = 16'h4675; w_imag[161] = 16'h9524;
w_real[162] = 16'h45CD; w_imag[162] = 16'h94B6;
w_real[163] = 16'h4524; w_imag[163] = 16'h9448;
w_real[164] = 16'h447A; w_imag[164] = 16'h93DC;
w_real[165] = 16'h43D0; w_imag[165] = 16'h9371;
w_real[166] = 16'h4325; w_imag[166] = 16'h9307;
w_real[167] = 16'h427A; w_imag[167] = 16'h929E;
w_real[168] = 16'h41CE; w_imag[168] = 16'h9236;
w_real[169] = 16'h4121; w_imag[169] = 16'h91D0;
w_real[170] = 16'h4073; w_imag[170] = 16'h916A;
w_real[171] = 16'h3FC5; w_imag[171] = 16'h9105;
w_real[172] = 16'h3F17; w_imag[172] = 16'h90A1;
w_real[173] = 16'h3E68; w_imag[173] = 16'h903F;
w_real[174] = 16'h3DB8; w_imag[174] = 16'h8FDD;
w_real[175] = 16'h3D07; w_imag[175] = 16'h8F7D;
w_real[176] = 16'h3C56; w_imag[176] = 16'h8F1E;
w_real[177] = 16'h3BA5; w_imag[177] = 16'h8EBF;
w_real[178] = 16'h3AF2; w_imag[178] = 16'h8E62;
w_real[179] = 16'h3A40; w_imag[179] = 16'h8E06;
w_real[180] = 16'h398C; w_imag[180] = 16'h8DAB;
w_real[181] = 16'h38D8; w_imag[181] = 16'h8D51;
w_real[182] = 16'h3824; w_imag[182] = 16'h8CF9;
w_real[183] = 16'h376F; w_imag[183] = 16'h8CA1;
w_real[184] = 16'h36BA; w_imag[184] = 16'h8C4B;
w_real[185] = 16'h3604; w_imag[185] = 16'h8BF5;
w_real[186] = 16'h354D; w_imag[186] = 16'h8BA1;
w_real[187] = 16'h3496; w_imag[187] = 16'h8B4E;
w_real[188] = 16'h33DE; w_imag[188] = 16'h8AFC;
w_real[189] = 16'h3326; w_imag[189] = 16'h8AAB;
w_real[190] = 16'h326E; w_imag[190] = 16'h8A5B;
w_real[191] = 16'h31B5; w_imag[191] = 16'h8A0C;
w_real[192] = 16'h30FB; w_imag[192] = 16'h89BF;
w_real[193] = 16'h3041; w_imag[193] = 16'h8972;
w_real[194] = 16'h2F87; w_imag[194] = 16'h8927;
w_real[195] = 16'h2ECC; w_imag[195] = 16'h88DD;
w_real[196] = 16'h2E11; w_imag[196] = 16'h8894;
w_real[197] = 16'h2D55; w_imag[197] = 16'h884C;
w_real[198] = 16'h2C98; w_imag[198] = 16'h8806;
w_real[199] = 16'h2BDC; w_imag[199] = 16'h87C0;
w_real[200] = 16'h2B1F; w_imag[200] = 16'h877C;
w_real[201] = 16'h2A61; w_imag[201] = 16'h8739;
w_real[202] = 16'h29A3; w_imag[202] = 16'h86F7;
w_real[203] = 16'h28E5; w_imag[203] = 16'h86B6;
w_real[204] = 16'h2826; w_imag[204] = 16'h8676;
w_real[205] = 16'h2767; w_imag[205] = 16'h8638;
w_real[206] = 16'h26A8; w_imag[206] = 16'h85FB;
w_real[207] = 16'h25E8; w_imag[207] = 16'h85BE;
w_real[208] = 16'h2528; w_imag[208] = 16'h8583;
w_real[209] = 16'h2467; w_imag[209] = 16'h854A;
w_real[210] = 16'h23A6; w_imag[210] = 16'h8511;
w_real[211] = 16'h22E5; w_imag[211] = 16'h84DA;
w_real[212] = 16'h2223; w_imag[212] = 16'h84A3;
w_real[213] = 16'h2161; w_imag[213] = 16'h846E;
w_real[214] = 16'h209F; w_imag[214] = 16'h843B;
w_real[215] = 16'h1FDC; w_imag[215] = 16'h8408;
w_real[216] = 16'h1F19; w_imag[216] = 16'h83D7;
w_real[217] = 16'h1E56; w_imag[217] = 16'h83A6;
w_real[218] = 16'h1D93; w_imag[218] = 16'h8377;
w_real[219] = 16'h1CCF; w_imag[219] = 16'h8349;
w_real[220] = 16'h1C0B; w_imag[220] = 16'h831D;
w_real[221] = 16'h1B47; w_imag[221] = 16'h82F1;
w_real[222] = 16'h1A82; w_imag[222] = 16'h82C7;
w_real[223] = 16'h19BD; w_imag[223] = 16'h829E;
w_real[224] = 16'h18F8; w_imag[224] = 16'h8276;
w_real[225] = 16'h1833; w_imag[225] = 16'h8250;
w_real[226] = 16'h176D; w_imag[226] = 16'h822A;
w_real[227] = 16'h16A8; w_imag[227] = 16'h8206;
w_real[228] = 16'h15E2; w_imag[228] = 16'h81E3;
w_real[229] = 16'h151B; w_imag[229] = 16'h81C1;
w_real[230] = 16'h1455; w_imag[230] = 16'h81A1;
w_real[231] = 16'h138E; w_imag[231] = 16'h8181;
w_real[232] = 16'h12C8; w_imag[232] = 16'h8163;
w_real[233] = 16'h1201; w_imag[233] = 16'h8146;
w_real[234] = 16'h1139; w_imag[234] = 16'h812B;
w_real[235] = 16'h1072; w_imag[235] = 16'h8110;
w_real[236] = 16'h0FAB; w_imag[236] = 16'h80F7;
w_real[237] = 16'h0EE3; w_imag[237] = 16'h80DF;
w_real[238] = 16'h0E1B; w_imag[238] = 16'h80C8;
w_real[239] = 16'h0D53; w_imag[239] = 16'h80B3;
w_real[240] = 16'h0C8B; w_imag[240] = 16'h809E;
w_real[241] = 16'h0BC3; w_imag[241] = 16'h808B;
w_real[242] = 16'h0AFB; w_imag[242] = 16'h8079;
w_real[243] = 16'h0A33; w_imag[243] = 16'h8069;
w_real[244] = 16'h096A; w_imag[244] = 16'h8059;
w_real[245] = 16'h08A2; w_imag[245] = 16'h804B;
w_real[246] = 16'h07D9; w_imag[246] = 16'h803E;
w_real[247] = 16'h0710; w_imag[247] = 16'h8032;
w_real[248] = 16'h0647; w_imag[248] = 16'h8028;
w_real[249] = 16'h057F; w_imag[249] = 16'h801F;
w_real[250] = 16'h04B6; w_imag[250] = 16'h8017;
w_real[251] = 16'h03ED; w_imag[251] = 16'h8010;
w_real[252] = 16'h0324; w_imag[252] = 16'h800A;
w_real[253] = 16'h025B; w_imag[253] = 16'h8006;
w_real[254] = 16'h0192; w_imag[254] = 16'h8003;
w_real[255] = 16'h00C9; w_imag[255] = 16'h8001;
w_real[256] = 16'h0000; w_imag[256] = 16'h8000;
w_real[257] = 16'hFF37; w_imag[257] = 16'h8001;
w_real[258] = 16'hFE6E; w_imag[258] = 16'h8003;
w_real[259] = 16'hFDA5; w_imag[259] = 16'h8006;
w_real[260] = 16'hFCDC; w_imag[260] = 16'h800A;
w_real[261] = 16'hFC13; w_imag[261] = 16'h8010;
w_real[262] = 16'hFB4A; w_imag[262] = 16'h8017;
w_real[263] = 16'hFA81; w_imag[263] = 16'h801F;
w_real[264] = 16'hF9B9; w_imag[264] = 16'h8028;
w_real[265] = 16'hF8F0; w_imag[265] = 16'h8032;
w_real[266] = 16'hF827; w_imag[266] = 16'h803E;
w_real[267] = 16'hF75E; w_imag[267] = 16'h804B;
w_real[268] = 16'hF696; w_imag[268] = 16'h8059;
w_real[269] = 16'hF5CD; w_imag[269] = 16'h8069;
w_real[270] = 16'hF505; w_imag[270] = 16'h8079;
w_real[271] = 16'hF43D; w_imag[271] = 16'h808B;
w_real[272] = 16'hF375; w_imag[272] = 16'h809E;
w_real[273] = 16'hF2AD; w_imag[273] = 16'h80B3;
w_real[274] = 16'hF1E5; w_imag[274] = 16'h80C8;
w_real[275] = 16'hF11D; w_imag[275] = 16'h80DF;
w_real[276] = 16'hF055; w_imag[276] = 16'h80F7;
w_real[277] = 16'hEF8E; w_imag[277] = 16'h8110;
w_real[278] = 16'hEEC7; w_imag[278] = 16'h812B;
w_real[279] = 16'hEDFF; w_imag[279] = 16'h8146;
w_real[280] = 16'hED38; w_imag[280] = 16'h8163;
w_real[281] = 16'hEC72; w_imag[281] = 16'h8181;
w_real[282] = 16'hEBAB; w_imag[282] = 16'h81A1;
w_real[283] = 16'hEAE5; w_imag[283] = 16'h81C1;
w_real[284] = 16'hEA1E; w_imag[284] = 16'h81E3;
w_real[285] = 16'hE958; w_imag[285] = 16'h8206;
w_real[286] = 16'hE893; w_imag[286] = 16'h822A;
w_real[287] = 16'hE7CD; w_imag[287] = 16'h8250;
w_real[288] = 16'hE708; w_imag[288] = 16'h8276;
w_real[289] = 16'hE643; w_imag[289] = 16'h829E;
w_real[290] = 16'hE57E; w_imag[290] = 16'h82C7;
w_real[291] = 16'hE4B9; w_imag[291] = 16'h82F1;
w_real[292] = 16'hE3F5; w_imag[292] = 16'h831D;
w_real[293] = 16'hE331; w_imag[293] = 16'h8349;
w_real[294] = 16'hE26D; w_imag[294] = 16'h8377;
w_real[295] = 16'hE1AA; w_imag[295] = 16'h83A6;
w_real[296] = 16'hE0E7; w_imag[296] = 16'h83D7;
w_real[297] = 16'hE024; w_imag[297] = 16'h8408;
w_real[298] = 16'hDF61; w_imag[298] = 16'h843B;
w_real[299] = 16'hDE9F; w_imag[299] = 16'h846E;
w_real[300] = 16'hDDDD; w_imag[300] = 16'h84A3;
w_real[301] = 16'hDD1B; w_imag[301] = 16'h84DA;
w_real[302] = 16'hDC5A; w_imag[302] = 16'h8511;
w_real[303] = 16'hDB99; w_imag[303] = 16'h854A;
w_real[304] = 16'hDAD8; w_imag[304] = 16'h8583;
w_real[305] = 16'hDA18; w_imag[305] = 16'h85BE;
w_real[306] = 16'hD958; w_imag[306] = 16'h85FB;
w_real[307] = 16'hD899; w_imag[307] = 16'h8638;
w_real[308] = 16'hD7DA; w_imag[308] = 16'h8676;
w_real[309] = 16'hD71B; w_imag[309] = 16'h86B6;
w_real[310] = 16'hD65D; w_imag[310] = 16'h86F7;
w_real[311] = 16'hD59F; w_imag[311] = 16'h8739;
w_real[312] = 16'hD4E1; w_imag[312] = 16'h877C;
w_real[313] = 16'hD424; w_imag[313] = 16'h87C0;
w_real[314] = 16'hD368; w_imag[314] = 16'h8806;
w_real[315] = 16'hD2AB; w_imag[315] = 16'h884C;
w_real[316] = 16'hD1EF; w_imag[316] = 16'h8894;
w_real[317] = 16'hD134; w_imag[317] = 16'h88DD;
w_real[318] = 16'hD079; w_imag[318] = 16'h8927;
w_real[319] = 16'hCFBF; w_imag[319] = 16'h8972;
w_real[320] = 16'hCF05; w_imag[320] = 16'h89BF;
w_real[321] = 16'hCE4B; w_imag[321] = 16'h8A0C;
w_real[322] = 16'hCD92; w_imag[322] = 16'h8A5B;
w_real[323] = 16'hCCDA; w_imag[323] = 16'h8AAB;
w_real[324] = 16'hCC22; w_imag[324] = 16'h8AFC;
w_real[325] = 16'hCB6A; w_imag[325] = 16'h8B4E;
w_real[326] = 16'hCAB3; w_imag[326] = 16'h8BA1;
w_real[327] = 16'hC9FC; w_imag[327] = 16'h8BF5;
w_real[328] = 16'hC946; w_imag[328] = 16'h8C4B;
w_real[329] = 16'hC891; w_imag[329] = 16'h8CA1;
w_real[330] = 16'hC7DC; w_imag[330] = 16'h8CF9;
w_real[331] = 16'hC728; w_imag[331] = 16'h8D51;
w_real[332] = 16'hC674; w_imag[332] = 16'h8DAB;
w_real[333] = 16'hC5C0; w_imag[333] = 16'h8E06;
w_real[334] = 16'hC50E; w_imag[334] = 16'h8E62;
w_real[335] = 16'hC45B; w_imag[335] = 16'h8EBF;
w_real[336] = 16'hC3AA; w_imag[336] = 16'h8F1E;
w_real[337] = 16'hC2F9; w_imag[337] = 16'h8F7D;
w_real[338] = 16'hC248; w_imag[338] = 16'h8FDD;
w_real[339] = 16'hC198; w_imag[339] = 16'h903F;
w_real[340] = 16'hC0E9; w_imag[340] = 16'h90A1;
w_real[341] = 16'hC03B; w_imag[341] = 16'h9105;
w_real[342] = 16'hBF8D; w_imag[342] = 16'h916A;
w_real[343] = 16'hBEDF; w_imag[343] = 16'h91D0;
w_real[344] = 16'hBE32; w_imag[344] = 16'h9236;
w_real[345] = 16'hBD86; w_imag[345] = 16'h929E;
w_real[346] = 16'hBCDB; w_imag[346] = 16'h9307;
w_real[347] = 16'hBC30; w_imag[347] = 16'h9371;
w_real[348] = 16'hBB86; w_imag[348] = 16'h93DC;
w_real[349] = 16'hBADC; w_imag[349] = 16'h9448;
w_real[350] = 16'hBA33; w_imag[350] = 16'h94B6;
w_real[351] = 16'hB98B; w_imag[351] = 16'h9524;
w_real[352] = 16'hB8E4; w_imag[352] = 16'h9593;
w_real[353] = 16'hB83D; w_imag[353] = 16'h9603;
w_real[354] = 16'hB797; w_imag[354] = 16'h9674;
w_real[355] = 16'hB6F1; w_imag[355] = 16'h96E7;
w_real[356] = 16'hB64C; w_imag[356] = 16'h975A;
w_real[357] = 16'hB5A8; w_imag[357] = 16'h97CE;
w_real[358] = 16'hB505; w_imag[358] = 16'h9843;
w_real[359] = 16'hB462; w_imag[359] = 16'h98BA;
w_real[360] = 16'hB3C1; w_imag[360] = 16'h9931;
w_real[361] = 16'hB31F; w_imag[361] = 16'h99A9;
w_real[362] = 16'hB27F; w_imag[362] = 16'h9A23;
w_real[363] = 16'hB1DF; w_imag[363] = 16'h9A9D;
w_real[364] = 16'hB141; w_imag[364] = 16'h9B18;
w_real[365] = 16'hB0A2; w_imag[365] = 16'h9B94;
w_real[366] = 16'hB005; w_imag[366] = 16'h9C11;
w_real[367] = 16'hAF69; w_imag[367] = 16'h9C8F;
w_real[368] = 16'hAECD; w_imag[368] = 16'h9D0E;
w_real[369] = 16'hAE32; w_imag[369] = 16'h9D8F;
w_real[370] = 16'hAD97; w_imag[370] = 16'h9E0F;
w_real[371] = 16'hACFE; w_imag[371] = 16'h9E91;
w_real[372] = 16'hAC65; w_imag[372] = 16'h9F14;
w_real[373] = 16'hABCD; w_imag[373] = 16'h9F98;
w_real[374] = 16'hAB36; w_imag[374] = 16'hA01D;
w_real[375] = 16'hAAA0; w_imag[375] = 16'hA0A2;
w_real[376] = 16'hAA0B; w_imag[376] = 16'hA129;
w_real[377] = 16'hA976; w_imag[377] = 16'hA1B0;
w_real[378] = 16'hA8E3; w_imag[378] = 16'hA239;
w_real[379] = 16'hA850; w_imag[379] = 16'hA2C2;
w_real[380] = 16'hA7BE; w_imag[380] = 16'hA34C;
w_real[381] = 16'hA72C; w_imag[381] = 16'hA3D7;
w_real[382] = 16'hA69C; w_imag[382] = 16'hA463;
w_real[383] = 16'hA60D; w_imag[383] = 16'hA4F0;
w_real[384] = 16'hA57E; w_imag[384] = 16'hA57E;
w_real[385] = 16'hA4F0; w_imag[385] = 16'hA60D;
w_real[386] = 16'hA463; w_imag[386] = 16'hA69C;
w_real[387] = 16'hA3D7; w_imag[387] = 16'hA72C;
w_real[388] = 16'hA34C; w_imag[388] = 16'hA7BE;
w_real[389] = 16'hA2C2; w_imag[389] = 16'hA850;
w_real[390] = 16'hA239; w_imag[390] = 16'hA8E3;
w_real[391] = 16'hA1B0; w_imag[391] = 16'hA976;
w_real[392] = 16'hA129; w_imag[392] = 16'hAA0B;
w_real[393] = 16'hA0A2; w_imag[393] = 16'hAAA0;
w_real[394] = 16'hA01D; w_imag[394] = 16'hAB36;
w_real[395] = 16'h9F98; w_imag[395] = 16'hABCD;
w_real[396] = 16'h9F14; w_imag[396] = 16'hAC65;
w_real[397] = 16'h9E91; w_imag[397] = 16'hACFE;
w_real[398] = 16'h9E0F; w_imag[398] = 16'hAD97;
w_real[399] = 16'h9D8F; w_imag[399] = 16'hAE32;
w_real[400] = 16'h9D0E; w_imag[400] = 16'hAECD;
w_real[401] = 16'h9C8F; w_imag[401] = 16'hAF69;
w_real[402] = 16'h9C11; w_imag[402] = 16'hB005;
w_real[403] = 16'h9B94; w_imag[403] = 16'hB0A2;
w_real[404] = 16'h9B18; w_imag[404] = 16'hB141;
w_real[405] = 16'h9A9D; w_imag[405] = 16'hB1DF;
w_real[406] = 16'h9A23; w_imag[406] = 16'hB27F;
w_real[407] = 16'h99A9; w_imag[407] = 16'hB31F;
w_real[408] = 16'h9931; w_imag[408] = 16'hB3C1;
w_real[409] = 16'h98BA; w_imag[409] = 16'hB462;
w_real[410] = 16'h9843; w_imag[410] = 16'hB505;
w_real[411] = 16'h97CE; w_imag[411] = 16'hB5A8;
w_real[412] = 16'h975A; w_imag[412] = 16'hB64C;
w_real[413] = 16'h96E7; w_imag[413] = 16'hB6F1;
w_real[414] = 16'h9674; w_imag[414] = 16'hB797;
w_real[415] = 16'h9603; w_imag[415] = 16'hB83D;
w_real[416] = 16'h9593; w_imag[416] = 16'hB8E4;
w_real[417] = 16'h9524; w_imag[417] = 16'hB98B;
w_real[418] = 16'h94B6; w_imag[418] = 16'hBA33;
w_real[419] = 16'h9448; w_imag[419] = 16'hBADC;
w_real[420] = 16'h93DC; w_imag[420] = 16'hBB86;
w_real[421] = 16'h9371; w_imag[421] = 16'hBC30;
w_real[422] = 16'h9307; w_imag[422] = 16'hBCDB;
w_real[423] = 16'h929E; w_imag[423] = 16'hBD86;
w_real[424] = 16'h9236; w_imag[424] = 16'hBE32;
w_real[425] = 16'h91D0; w_imag[425] = 16'hBEDF;
w_real[426] = 16'h916A; w_imag[426] = 16'hBF8D;
w_real[427] = 16'h9105; w_imag[427] = 16'hC03B;
w_real[428] = 16'h90A1; w_imag[428] = 16'hC0E9;
w_real[429] = 16'h903F; w_imag[429] = 16'hC198;
w_real[430] = 16'h8FDD; w_imag[430] = 16'hC248;
w_real[431] = 16'h8F7D; w_imag[431] = 16'hC2F9;
w_real[432] = 16'h8F1E; w_imag[432] = 16'hC3AA;
w_real[433] = 16'h8EBF; w_imag[433] = 16'hC45B;
w_real[434] = 16'h8E62; w_imag[434] = 16'hC50E;
w_real[435] = 16'h8E06; w_imag[435] = 16'hC5C0;
w_real[436] = 16'h8DAB; w_imag[436] = 16'hC674;
w_real[437] = 16'h8D51; w_imag[437] = 16'hC728;
w_real[438] = 16'h8CF9; w_imag[438] = 16'hC7DC;
w_real[439] = 16'h8CA1; w_imag[439] = 16'hC891;
w_real[440] = 16'h8C4B; w_imag[440] = 16'hC946;
w_real[441] = 16'h8BF5; w_imag[441] = 16'hC9FC;
w_real[442] = 16'h8BA1; w_imag[442] = 16'hCAB3;
w_real[443] = 16'h8B4E; w_imag[443] = 16'hCB6A;
w_real[444] = 16'h8AFC; w_imag[444] = 16'hCC22;
w_real[445] = 16'h8AAB; w_imag[445] = 16'hCCDA;
w_real[446] = 16'h8A5B; w_imag[446] = 16'hCD92;
w_real[447] = 16'h8A0C; w_imag[447] = 16'hCE4B;
w_real[448] = 16'h89BF; w_imag[448] = 16'hCF05;
w_real[449] = 16'h8972; w_imag[449] = 16'hCFBF;
w_real[450] = 16'h8927; w_imag[450] = 16'hD079;
w_real[451] = 16'h88DD; w_imag[451] = 16'hD134;
w_real[452] = 16'h8894; w_imag[452] = 16'hD1EF;
w_real[453] = 16'h884C; w_imag[453] = 16'hD2AB;
w_real[454] = 16'h8806; w_imag[454] = 16'hD368;
w_real[455] = 16'h87C0; w_imag[455] = 16'hD424;
w_real[456] = 16'h877C; w_imag[456] = 16'hD4E1;
w_real[457] = 16'h8739; w_imag[457] = 16'hD59F;
w_real[458] = 16'h86F7; w_imag[458] = 16'hD65D;
w_real[459] = 16'h86B6; w_imag[459] = 16'hD71B;
w_real[460] = 16'h8676; w_imag[460] = 16'hD7DA;
w_real[461] = 16'h8638; w_imag[461] = 16'hD899;
w_real[462] = 16'h85FB; w_imag[462] = 16'hD958;
w_real[463] = 16'h85BE; w_imag[463] = 16'hDA18;
w_real[464] = 16'h8583; w_imag[464] = 16'hDAD8;
w_real[465] = 16'h854A; w_imag[465] = 16'hDB99;
w_real[466] = 16'h8511; w_imag[466] = 16'hDC5A;
w_real[467] = 16'h84DA; w_imag[467] = 16'hDD1B;
w_real[468] = 16'h84A3; w_imag[468] = 16'hDDDD;
w_real[469] = 16'h846E; w_imag[469] = 16'hDE9F;
w_real[470] = 16'h843B; w_imag[470] = 16'hDF61;
w_real[471] = 16'h8408; w_imag[471] = 16'hE024;
w_real[472] = 16'h83D7; w_imag[472] = 16'hE0E7;
w_real[473] = 16'h83A6; w_imag[473] = 16'hE1AA;
w_real[474] = 16'h8377; w_imag[474] = 16'hE26D;
w_real[475] = 16'h8349; w_imag[475] = 16'hE331;
w_real[476] = 16'h831D; w_imag[476] = 16'hE3F5;
w_real[477] = 16'h82F1; w_imag[477] = 16'hE4B9;
w_real[478] = 16'h82C7; w_imag[478] = 16'hE57E;
w_real[479] = 16'h829E; w_imag[479] = 16'hE643;
w_real[480] = 16'h8276; w_imag[480] = 16'hE708;
w_real[481] = 16'h8250; w_imag[481] = 16'hE7CD;
w_real[482] = 16'h822A; w_imag[482] = 16'hE893;
w_real[483] = 16'h8206; w_imag[483] = 16'hE958;
w_real[484] = 16'h81E3; w_imag[484] = 16'hEA1E;
w_real[485] = 16'h81C1; w_imag[485] = 16'hEAE5;
w_real[486] = 16'h81A1; w_imag[486] = 16'hEBAB;
w_real[487] = 16'h8181; w_imag[487] = 16'hEC72;
w_real[488] = 16'h8163; w_imag[488] = 16'hED38;
w_real[489] = 16'h8146; w_imag[489] = 16'hEDFF;
w_real[490] = 16'h812B; w_imag[490] = 16'hEEC7;
w_real[491] = 16'h8110; w_imag[491] = 16'hEF8E;
w_real[492] = 16'h80F7; w_imag[492] = 16'hF055;
w_real[493] = 16'h80DF; w_imag[493] = 16'hF11D;
w_real[494] = 16'h80C8; w_imag[494] = 16'hF1E5;
w_real[495] = 16'h80B3; w_imag[495] = 16'hF2AD;
w_real[496] = 16'h809E; w_imag[496] = 16'hF375;
w_real[497] = 16'h808B; w_imag[497] = 16'hF43D;
w_real[498] = 16'h8079; w_imag[498] = 16'hF505;
w_real[499] = 16'h8069; w_imag[499] = 16'hF5CD;
w_real[500] = 16'h8059; w_imag[500] = 16'hF696;
w_real[501] = 16'h804B; w_imag[501] = 16'hF75E;
w_real[502] = 16'h803E; w_imag[502] = 16'hF827;
w_real[503] = 16'h8032; w_imag[503] = 16'hF8F0;
w_real[504] = 16'h8028; w_imag[504] = 16'hF9B9;
w_real[505] = 16'h801F; w_imag[505] = 16'hFA81;
w_real[506] = 16'h8017; w_imag[506] = 16'hFB4A;
w_real[507] = 16'h8010; w_imag[507] = 16'hFC13;
w_real[508] = 16'h800A; w_imag[508] = 16'hFCDC;
w_real[509] = 16'h8006; w_imag[509] = 16'hFDA5;
w_real[510] = 16'h8003; w_imag[510] = 16'hFE6E;
w_real[511] = 16'h8001; w_imag[511] = 16'hFF37;
w_real[512] = 16'h8000; w_imag[512] = 16'h0000;
w_real[513] = 16'h8001; w_imag[513] = 16'h00C9;
w_real[514] = 16'h8003; w_imag[514] = 16'h0192;
w_real[515] = 16'h8006; w_imag[515] = 16'h025B;
w_real[516] = 16'h800A; w_imag[516] = 16'h0324;
w_real[517] = 16'h8010; w_imag[517] = 16'h03ED;
w_real[518] = 16'h8017; w_imag[518] = 16'h04B6;
w_real[519] = 16'h801F; w_imag[519] = 16'h057F;
w_real[520] = 16'h8028; w_imag[520] = 16'h0647;
w_real[521] = 16'h8032; w_imag[521] = 16'h0710;
w_real[522] = 16'h803E; w_imag[522] = 16'h07D9;
w_real[523] = 16'h804B; w_imag[523] = 16'h08A2;
w_real[524] = 16'h8059; w_imag[524] = 16'h096A;
w_real[525] = 16'h8069; w_imag[525] = 16'h0A33;
w_real[526] = 16'h8079; w_imag[526] = 16'h0AFB;
w_real[527] = 16'h808B; w_imag[527] = 16'h0BC3;
w_real[528] = 16'h809E; w_imag[528] = 16'h0C8B;
w_real[529] = 16'h80B3; w_imag[529] = 16'h0D53;
w_real[530] = 16'h80C8; w_imag[530] = 16'h0E1B;
w_real[531] = 16'h80DF; w_imag[531] = 16'h0EE3;
w_real[532] = 16'h80F7; w_imag[532] = 16'h0FAB;
w_real[533] = 16'h8110; w_imag[533] = 16'h1072;
w_real[534] = 16'h812B; w_imag[534] = 16'h1139;
w_real[535] = 16'h8146; w_imag[535] = 16'h1201;
w_real[536] = 16'h8163; w_imag[536] = 16'h12C8;
w_real[537] = 16'h8181; w_imag[537] = 16'h138E;
w_real[538] = 16'h81A1; w_imag[538] = 16'h1455;
w_real[539] = 16'h81C1; w_imag[539] = 16'h151B;
w_real[540] = 16'h81E3; w_imag[540] = 16'h15E2;
w_real[541] = 16'h8206; w_imag[541] = 16'h16A8;
w_real[542] = 16'h822A; w_imag[542] = 16'h176D;
w_real[543] = 16'h8250; w_imag[543] = 16'h1833;
w_real[544] = 16'h8276; w_imag[544] = 16'h18F8;
w_real[545] = 16'h829E; w_imag[545] = 16'h19BD;
w_real[546] = 16'h82C7; w_imag[546] = 16'h1A82;
w_real[547] = 16'h82F1; w_imag[547] = 16'h1B47;
w_real[548] = 16'h831D; w_imag[548] = 16'h1C0B;
w_real[549] = 16'h8349; w_imag[549] = 16'h1CCF;
w_real[550] = 16'h8377; w_imag[550] = 16'h1D93;
w_real[551] = 16'h83A6; w_imag[551] = 16'h1E56;
w_real[552] = 16'h83D7; w_imag[552] = 16'h1F19;
w_real[553] = 16'h8408; w_imag[553] = 16'h1FDC;
w_real[554] = 16'h843B; w_imag[554] = 16'h209F;
w_real[555] = 16'h846E; w_imag[555] = 16'h2161;
w_real[556] = 16'h84A3; w_imag[556] = 16'h2223;
w_real[557] = 16'h84DA; w_imag[557] = 16'h22E5;
w_real[558] = 16'h8511; w_imag[558] = 16'h23A6;
w_real[559] = 16'h854A; w_imag[559] = 16'h2467;
w_real[560] = 16'h8583; w_imag[560] = 16'h2528;
w_real[561] = 16'h85BE; w_imag[561] = 16'h25E8;
w_real[562] = 16'h85FB; w_imag[562] = 16'h26A8;
w_real[563] = 16'h8638; w_imag[563] = 16'h2767;
w_real[564] = 16'h8676; w_imag[564] = 16'h2826;
w_real[565] = 16'h86B6; w_imag[565] = 16'h28E5;
w_real[566] = 16'h86F7; w_imag[566] = 16'h29A3;
w_real[567] = 16'h8739; w_imag[567] = 16'h2A61;
w_real[568] = 16'h877C; w_imag[568] = 16'h2B1F;
w_real[569] = 16'h87C0; w_imag[569] = 16'h2BDC;
w_real[570] = 16'h8806; w_imag[570] = 16'h2C98;
w_real[571] = 16'h884C; w_imag[571] = 16'h2D55;
w_real[572] = 16'h8894; w_imag[572] = 16'h2E11;
w_real[573] = 16'h88DD; w_imag[573] = 16'h2ECC;
w_real[574] = 16'h8927; w_imag[574] = 16'h2F87;
w_real[575] = 16'h8972; w_imag[575] = 16'h3041;
w_real[576] = 16'h89BF; w_imag[576] = 16'h30FB;
w_real[577] = 16'h8A0C; w_imag[577] = 16'h31B5;
w_real[578] = 16'h8A5B; w_imag[578] = 16'h326E;
w_real[579] = 16'h8AAB; w_imag[579] = 16'h3326;
w_real[580] = 16'h8AFC; w_imag[580] = 16'h33DE;
w_real[581] = 16'h8B4E; w_imag[581] = 16'h3496;
w_real[582] = 16'h8BA1; w_imag[582] = 16'h354D;
w_real[583] = 16'h8BF5; w_imag[583] = 16'h3604;
w_real[584] = 16'h8C4B; w_imag[584] = 16'h36BA;
w_real[585] = 16'h8CA1; w_imag[585] = 16'h376F;
w_real[586] = 16'h8CF9; w_imag[586] = 16'h3824;
w_real[587] = 16'h8D51; w_imag[587] = 16'h38D8;
w_real[588] = 16'h8DAB; w_imag[588] = 16'h398C;
w_real[589] = 16'h8E06; w_imag[589] = 16'h3A40;
w_real[590] = 16'h8E62; w_imag[590] = 16'h3AF2;
w_real[591] = 16'h8EBF; w_imag[591] = 16'h3BA5;
w_real[592] = 16'h8F1E; w_imag[592] = 16'h3C56;
w_real[593] = 16'h8F7D; w_imag[593] = 16'h3D07;
w_real[594] = 16'h8FDD; w_imag[594] = 16'h3DB8;
w_real[595] = 16'h903F; w_imag[595] = 16'h3E68;
w_real[596] = 16'h90A1; w_imag[596] = 16'h3F17;
w_real[597] = 16'h9105; w_imag[597] = 16'h3FC5;
w_real[598] = 16'h916A; w_imag[598] = 16'h4073;
w_real[599] = 16'h91D0; w_imag[599] = 16'h4121;
w_real[600] = 16'h9236; w_imag[600] = 16'h41CE;
w_real[601] = 16'h929E; w_imag[601] = 16'h427A;
w_real[602] = 16'h9307; w_imag[602] = 16'h4325;
w_real[603] = 16'h9371; w_imag[603] = 16'h43D0;
w_real[604] = 16'h93DC; w_imag[604] = 16'h447A;
w_real[605] = 16'h9448; w_imag[605] = 16'h4524;
w_real[606] = 16'h94B6; w_imag[606] = 16'h45CD;
w_real[607] = 16'h9524; w_imag[607] = 16'h4675;
w_real[608] = 16'h9593; w_imag[608] = 16'h471C;
w_real[609] = 16'h9603; w_imag[609] = 16'h47C3;
w_real[610] = 16'h9674; w_imag[610] = 16'h4869;
w_real[611] = 16'h96E7; w_imag[611] = 16'h490F;
w_real[612] = 16'h975A; w_imag[612] = 16'h49B4;
w_real[613] = 16'h97CE; w_imag[613] = 16'h4A58;
w_real[614] = 16'h9843; w_imag[614] = 16'h4AFB;
w_real[615] = 16'h98BA; w_imag[615] = 16'h4B9E;
w_real[616] = 16'h9931; w_imag[616] = 16'h4C3F;
w_real[617] = 16'h99A9; w_imag[617] = 16'h4CE1;
w_real[618] = 16'h9A23; w_imag[618] = 16'h4D81;
w_real[619] = 16'h9A9D; w_imag[619] = 16'h4E21;
w_real[620] = 16'h9B18; w_imag[620] = 16'h4EBF;
w_real[621] = 16'h9B94; w_imag[621] = 16'h4F5E;
w_real[622] = 16'h9C11; w_imag[622] = 16'h4FFB;
w_real[623] = 16'h9C8F; w_imag[623] = 16'h5097;
w_real[624] = 16'h9D0E; w_imag[624] = 16'h5133;
w_real[625] = 16'h9D8F; w_imag[625] = 16'h51CE;
w_real[626] = 16'h9E0F; w_imag[626] = 16'h5269;
w_real[627] = 16'h9E91; w_imag[627] = 16'h5302;
w_real[628] = 16'h9F14; w_imag[628] = 16'h539B;
w_real[629] = 16'h9F98; w_imag[629] = 16'h5433;
w_real[630] = 16'hA01D; w_imag[630] = 16'h54CA;
w_real[631] = 16'hA0A2; w_imag[631] = 16'h5560;
w_real[632] = 16'hA129; w_imag[632] = 16'h55F5;
w_real[633] = 16'hA1B0; w_imag[633] = 16'h568A;
w_real[634] = 16'hA239; w_imag[634] = 16'h571D;
w_real[635] = 16'hA2C2; w_imag[635] = 16'h57B0;
w_real[636] = 16'hA34C; w_imag[636] = 16'h5842;
w_real[637] = 16'hA3D7; w_imag[637] = 16'h58D4;
w_real[638] = 16'hA463; w_imag[638] = 16'h5964;
w_real[639] = 16'hA4F0; w_imag[639] = 16'h59F3;
w_real[640] = 16'hA57E; w_imag[640] = 16'h5A82;
w_real[641] = 16'hA60D; w_imag[641] = 16'h5B10;
w_real[642] = 16'hA69C; w_imag[642] = 16'h5B9D;
w_real[643] = 16'hA72C; w_imag[643] = 16'h5C29;
w_real[644] = 16'hA7BE; w_imag[644] = 16'h5CB4;
w_real[645] = 16'hA850; w_imag[645] = 16'h5D3E;
w_real[646] = 16'hA8E3; w_imag[646] = 16'h5DC7;
w_real[647] = 16'hA976; w_imag[647] = 16'h5E50;
w_real[648] = 16'hAA0B; w_imag[648] = 16'h5ED7;
w_real[649] = 16'hAAA0; w_imag[649] = 16'h5F5E;
w_real[650] = 16'hAB36; w_imag[650] = 16'h5FE3;
w_real[651] = 16'hABCD; w_imag[651] = 16'h6068;
w_real[652] = 16'hAC65; w_imag[652] = 16'h60EC;
w_real[653] = 16'hACFE; w_imag[653] = 16'h616F;
w_real[654] = 16'hAD97; w_imag[654] = 16'h61F1;
w_real[655] = 16'hAE32; w_imag[655] = 16'h6271;
w_real[656] = 16'hAECD; w_imag[656] = 16'h62F2;
w_real[657] = 16'hAF69; w_imag[657] = 16'h6371;
w_real[658] = 16'hB005; w_imag[658] = 16'h63EF;
w_real[659] = 16'hB0A2; w_imag[659] = 16'h646C;
w_real[660] = 16'hB141; w_imag[660] = 16'h64E8;
w_real[661] = 16'hB1DF; w_imag[661] = 16'h6563;
w_real[662] = 16'hB27F; w_imag[662] = 16'h65DD;
w_real[663] = 16'hB31F; w_imag[663] = 16'h6657;
w_real[664] = 16'hB3C1; w_imag[664] = 16'h66CF;
w_real[665] = 16'hB462; w_imag[665] = 16'h6746;
w_real[666] = 16'hB505; w_imag[666] = 16'h67BD;
w_real[667] = 16'hB5A8; w_imag[667] = 16'h6832;
w_real[668] = 16'hB64C; w_imag[668] = 16'h68A6;
w_real[669] = 16'hB6F1; w_imag[669] = 16'h6919;
w_real[670] = 16'hB797; w_imag[670] = 16'h698C;
w_real[671] = 16'hB83D; w_imag[671] = 16'h69FD;
w_real[672] = 16'hB8E4; w_imag[672] = 16'h6A6D;
w_real[673] = 16'hB98B; w_imag[673] = 16'h6ADC;
w_real[674] = 16'hBA33; w_imag[674] = 16'h6B4A;
w_real[675] = 16'hBADC; w_imag[675] = 16'h6BB8;
w_real[676] = 16'hBB86; w_imag[676] = 16'h6C24;
w_real[677] = 16'hBC30; w_imag[677] = 16'h6C8F;
w_real[678] = 16'hBCDB; w_imag[678] = 16'h6CF9;
w_real[679] = 16'hBD86; w_imag[679] = 16'h6D62;
w_real[680] = 16'hBE32; w_imag[680] = 16'h6DCA;
w_real[681] = 16'hBEDF; w_imag[681] = 16'h6E30;
w_real[682] = 16'hBF8D; w_imag[682] = 16'h6E96;
w_real[683] = 16'hC03B; w_imag[683] = 16'h6EFB;
w_real[684] = 16'hC0E9; w_imag[684] = 16'h6F5F;
w_real[685] = 16'hC198; w_imag[685] = 16'h6FC1;
w_real[686] = 16'hC248; w_imag[686] = 16'h7023;
w_real[687] = 16'hC2F9; w_imag[687] = 16'h7083;
w_real[688] = 16'hC3AA; w_imag[688] = 16'h70E2;
w_real[689] = 16'hC45B; w_imag[689] = 16'h7141;
w_real[690] = 16'hC50E; w_imag[690] = 16'h719E;
w_real[691] = 16'hC5C0; w_imag[691] = 16'h71FA;
w_real[692] = 16'hC674; w_imag[692] = 16'h7255;
w_real[693] = 16'hC728; w_imag[693] = 16'h72AF;
w_real[694] = 16'hC7DC; w_imag[694] = 16'h7307;
w_real[695] = 16'hC891; w_imag[695] = 16'h735F;
w_real[696] = 16'hC946; w_imag[696] = 16'h73B5;
w_real[697] = 16'hC9FC; w_imag[697] = 16'h740B;
w_real[698] = 16'hCAB3; w_imag[698] = 16'h745F;
w_real[699] = 16'hCB6A; w_imag[699] = 16'h74B2;
w_real[700] = 16'hCC22; w_imag[700] = 16'h7504;
w_real[701] = 16'hCCDA; w_imag[701] = 16'h7555;
w_real[702] = 16'hCD92; w_imag[702] = 16'h75A5;
w_real[703] = 16'hCE4B; w_imag[703] = 16'h75F4;
w_real[704] = 16'hCF05; w_imag[704] = 16'h7641;
w_real[705] = 16'hCFBF; w_imag[705] = 16'h768E;
w_real[706] = 16'hD079; w_imag[706] = 16'h76D9;
w_real[707] = 16'hD134; w_imag[707] = 16'h7723;
w_real[708] = 16'hD1EF; w_imag[708] = 16'h776C;
w_real[709] = 16'hD2AB; w_imag[709] = 16'h77B4;
w_real[710] = 16'hD368; w_imag[710] = 16'h77FA;
w_real[711] = 16'hD424; w_imag[711] = 16'h7840;
w_real[712] = 16'hD4E1; w_imag[712] = 16'h7884;
w_real[713] = 16'hD59F; w_imag[713] = 16'h78C7;
w_real[714] = 16'hD65D; w_imag[714] = 16'h7909;
w_real[715] = 16'hD71B; w_imag[715] = 16'h794A;
w_real[716] = 16'hD7DA; w_imag[716] = 16'h798A;
w_real[717] = 16'hD899; w_imag[717] = 16'h79C8;
w_real[718] = 16'hD958; w_imag[718] = 16'h7A05;
w_real[719] = 16'hDA18; w_imag[719] = 16'h7A42;
w_real[720] = 16'hDAD8; w_imag[720] = 16'h7A7D;
w_real[721] = 16'hDB99; w_imag[721] = 16'h7AB6;
w_real[722] = 16'hDC5A; w_imag[722] = 16'h7AEF;
w_real[723] = 16'hDD1B; w_imag[723] = 16'h7B26;
w_real[724] = 16'hDDDD; w_imag[724] = 16'h7B5D;
w_real[725] = 16'hDE9F; w_imag[725] = 16'h7B92;
w_real[726] = 16'hDF61; w_imag[726] = 16'h7BC5;
w_real[727] = 16'hE024; w_imag[727] = 16'h7BF8;
w_real[728] = 16'hE0E7; w_imag[728] = 16'h7C29;
w_real[729] = 16'hE1AA; w_imag[729] = 16'h7C5A;
w_real[730] = 16'hE26D; w_imag[730] = 16'h7C89;
w_real[731] = 16'hE331; w_imag[731] = 16'h7CB7;
w_real[732] = 16'hE3F5; w_imag[732] = 16'h7CE3;
w_real[733] = 16'hE4B9; w_imag[733] = 16'h7D0F;
w_real[734] = 16'hE57E; w_imag[734] = 16'h7D39;
w_real[735] = 16'hE643; w_imag[735] = 16'h7D62;
w_real[736] = 16'hE708; w_imag[736] = 16'h7D8A;
w_real[737] = 16'hE7CD; w_imag[737] = 16'h7DB0;
w_real[738] = 16'hE893; w_imag[738] = 16'h7DD6;
w_real[739] = 16'hE958; w_imag[739] = 16'h7DFA;
w_real[740] = 16'hEA1E; w_imag[740] = 16'h7E1D;
w_real[741] = 16'hEAE5; w_imag[741] = 16'h7E3F;
w_real[742] = 16'hEBAB; w_imag[742] = 16'h7E5F;
w_real[743] = 16'hEC72; w_imag[743] = 16'h7E7F;
w_real[744] = 16'hED38; w_imag[744] = 16'h7E9D;
w_real[745] = 16'hEDFF; w_imag[745] = 16'h7EBA;
w_real[746] = 16'hEEC7; w_imag[746] = 16'h7ED5;
w_real[747] = 16'hEF8E; w_imag[747] = 16'h7EF0;
w_real[748] = 16'hF055; w_imag[748] = 16'h7F09;
w_real[749] = 16'hF11D; w_imag[749] = 16'h7F21;
w_real[750] = 16'hF1E5; w_imag[750] = 16'h7F38;
w_real[751] = 16'hF2AD; w_imag[751] = 16'h7F4D;
w_real[752] = 16'hF375; w_imag[752] = 16'h7F62;
w_real[753] = 16'hF43D; w_imag[753] = 16'h7F75;
w_real[754] = 16'hF505; w_imag[754] = 16'h7F87;
w_real[755] = 16'hF5CD; w_imag[755] = 16'h7F97;
w_real[756] = 16'hF696; w_imag[756] = 16'h7FA7;
w_real[757] = 16'hF75E; w_imag[757] = 16'h7FB5;
w_real[758] = 16'hF827; w_imag[758] = 16'h7FC2;
w_real[759] = 16'hF8F0; w_imag[759] = 16'h7FCE;
w_real[760] = 16'hF9B9; w_imag[760] = 16'h7FD8;
w_real[761] = 16'hFA81; w_imag[761] = 16'h7FE1;
w_real[762] = 16'hFB4A; w_imag[762] = 16'h7FE9;
w_real[763] = 16'hFC13; w_imag[763] = 16'h7FF0;
w_real[764] = 16'hFCDC; w_imag[764] = 16'h7FF6;
w_real[765] = 16'hFDA5; w_imag[765] = 16'h7FFA;
w_real[766] = 16'hFE6E; w_imag[766] = 16'h7FFD;
w_real[767] = 16'hFF37; w_imag[767] = 16'h7FFF;
w_real[768] = 16'h0000; w_imag[768] = 16'h7FFF;
w_real[769] = 16'h00C9; w_imag[769] = 16'h7FFF;
w_real[770] = 16'h0192; w_imag[770] = 16'h7FFD;
w_real[771] = 16'h025B; w_imag[771] = 16'h7FFA;
w_real[772] = 16'h0324; w_imag[772] = 16'h7FF6;
w_real[773] = 16'h03ED; w_imag[773] = 16'h7FF0;
w_real[774] = 16'h04B6; w_imag[774] = 16'h7FE9;
w_real[775] = 16'h057F; w_imag[775] = 16'h7FE1;
w_real[776] = 16'h0647; w_imag[776] = 16'h7FD8;
w_real[777] = 16'h0710; w_imag[777] = 16'h7FCE;
w_real[778] = 16'h07D9; w_imag[778] = 16'h7FC2;
w_real[779] = 16'h08A2; w_imag[779] = 16'h7FB5;
w_real[780] = 16'h096A; w_imag[780] = 16'h7FA7;
w_real[781] = 16'h0A33; w_imag[781] = 16'h7F97;
w_real[782] = 16'h0AFB; w_imag[782] = 16'h7F87;
w_real[783] = 16'h0BC3; w_imag[783] = 16'h7F75;
w_real[784] = 16'h0C8B; w_imag[784] = 16'h7F62;
w_real[785] = 16'h0D53; w_imag[785] = 16'h7F4D;
w_real[786] = 16'h0E1B; w_imag[786] = 16'h7F38;
w_real[787] = 16'h0EE3; w_imag[787] = 16'h7F21;
w_real[788] = 16'h0FAB; w_imag[788] = 16'h7F09;
w_real[789] = 16'h1072; w_imag[789] = 16'h7EF0;
w_real[790] = 16'h1139; w_imag[790] = 16'h7ED5;
w_real[791] = 16'h1201; w_imag[791] = 16'h7EBA;
w_real[792] = 16'h12C8; w_imag[792] = 16'h7E9D;
w_real[793] = 16'h138E; w_imag[793] = 16'h7E7F;
w_real[794] = 16'h1455; w_imag[794] = 16'h7E5F;
w_real[795] = 16'h151B; w_imag[795] = 16'h7E3F;
w_real[796] = 16'h15E2; w_imag[796] = 16'h7E1D;
w_real[797] = 16'h16A8; w_imag[797] = 16'h7DFA;
w_real[798] = 16'h176D; w_imag[798] = 16'h7DD6;
w_real[799] = 16'h1833; w_imag[799] = 16'h7DB0;
w_real[800] = 16'h18F8; w_imag[800] = 16'h7D8A;
w_real[801] = 16'h19BD; w_imag[801] = 16'h7D62;
w_real[802] = 16'h1A82; w_imag[802] = 16'h7D39;
w_real[803] = 16'h1B47; w_imag[803] = 16'h7D0F;
w_real[804] = 16'h1C0B; w_imag[804] = 16'h7CE3;
w_real[805] = 16'h1CCF; w_imag[805] = 16'h7CB7;
w_real[806] = 16'h1D93; w_imag[806] = 16'h7C89;
w_real[807] = 16'h1E56; w_imag[807] = 16'h7C5A;
w_real[808] = 16'h1F19; w_imag[808] = 16'h7C29;
w_real[809] = 16'h1FDC; w_imag[809] = 16'h7BF8;
w_real[810] = 16'h209F; w_imag[810] = 16'h7BC5;
w_real[811] = 16'h2161; w_imag[811] = 16'h7B92;
w_real[812] = 16'h2223; w_imag[812] = 16'h7B5D;
w_real[813] = 16'h22E5; w_imag[813] = 16'h7B26;
w_real[814] = 16'h23A6; w_imag[814] = 16'h7AEF;
w_real[815] = 16'h2467; w_imag[815] = 16'h7AB6;
w_real[816] = 16'h2528; w_imag[816] = 16'h7A7D;
w_real[817] = 16'h25E8; w_imag[817] = 16'h7A42;
w_real[818] = 16'h26A8; w_imag[818] = 16'h7A05;
w_real[819] = 16'h2767; w_imag[819] = 16'h79C8;
w_real[820] = 16'h2826; w_imag[820] = 16'h798A;
w_real[821] = 16'h28E5; w_imag[821] = 16'h794A;
w_real[822] = 16'h29A3; w_imag[822] = 16'h7909;
w_real[823] = 16'h2A61; w_imag[823] = 16'h78C7;
w_real[824] = 16'h2B1F; w_imag[824] = 16'h7884;
w_real[825] = 16'h2BDC; w_imag[825] = 16'h7840;
w_real[826] = 16'h2C98; w_imag[826] = 16'h77FA;
w_real[827] = 16'h2D55; w_imag[827] = 16'h77B4;
w_real[828] = 16'h2E11; w_imag[828] = 16'h776C;
w_real[829] = 16'h2ECC; w_imag[829] = 16'h7723;
w_real[830] = 16'h2F87; w_imag[830] = 16'h76D9;
w_real[831] = 16'h3041; w_imag[831] = 16'h768E;
w_real[832] = 16'h30FB; w_imag[832] = 16'h7641;
w_real[833] = 16'h31B5; w_imag[833] = 16'h75F4;
w_real[834] = 16'h326E; w_imag[834] = 16'h75A5;
w_real[835] = 16'h3326; w_imag[835] = 16'h7555;
w_real[836] = 16'h33DE; w_imag[836] = 16'h7504;
w_real[837] = 16'h3496; w_imag[837] = 16'h74B2;
w_real[838] = 16'h354D; w_imag[838] = 16'h745F;
w_real[839] = 16'h3604; w_imag[839] = 16'h740B;
w_real[840] = 16'h36BA; w_imag[840] = 16'h73B5;
w_real[841] = 16'h376F; w_imag[841] = 16'h735F;
w_real[842] = 16'h3824; w_imag[842] = 16'h7307;
w_real[843] = 16'h38D8; w_imag[843] = 16'h72AF;
w_real[844] = 16'h398C; w_imag[844] = 16'h7255;
w_real[845] = 16'h3A40; w_imag[845] = 16'h71FA;
w_real[846] = 16'h3AF2; w_imag[846] = 16'h719E;
w_real[847] = 16'h3BA5; w_imag[847] = 16'h7141;
w_real[848] = 16'h3C56; w_imag[848] = 16'h70E2;
w_real[849] = 16'h3D07; w_imag[849] = 16'h7083;
w_real[850] = 16'h3DB8; w_imag[850] = 16'h7023;
w_real[851] = 16'h3E68; w_imag[851] = 16'h6FC1;
w_real[852] = 16'h3F17; w_imag[852] = 16'h6F5F;
w_real[853] = 16'h3FC5; w_imag[853] = 16'h6EFB;
w_real[854] = 16'h4073; w_imag[854] = 16'h6E96;
w_real[855] = 16'h4121; w_imag[855] = 16'h6E30;
w_real[856] = 16'h41CE; w_imag[856] = 16'h6DCA;
w_real[857] = 16'h427A; w_imag[857] = 16'h6D62;
w_real[858] = 16'h4325; w_imag[858] = 16'h6CF9;
w_real[859] = 16'h43D0; w_imag[859] = 16'h6C8F;
w_real[860] = 16'h447A; w_imag[860] = 16'h6C24;
w_real[861] = 16'h4524; w_imag[861] = 16'h6BB8;
w_real[862] = 16'h45CD; w_imag[862] = 16'h6B4A;
w_real[863] = 16'h4675; w_imag[863] = 16'h6ADC;
w_real[864] = 16'h471C; w_imag[864] = 16'h6A6D;
w_real[865] = 16'h47C3; w_imag[865] = 16'h69FD;
w_real[866] = 16'h4869; w_imag[866] = 16'h698C;
w_real[867] = 16'h490F; w_imag[867] = 16'h6919;
w_real[868] = 16'h49B4; w_imag[868] = 16'h68A6;
w_real[869] = 16'h4A58; w_imag[869] = 16'h6832;
w_real[870] = 16'h4AFB; w_imag[870] = 16'h67BD;
w_real[871] = 16'h4B9E; w_imag[871] = 16'h6746;
w_real[872] = 16'h4C3F; w_imag[872] = 16'h66CF;
w_real[873] = 16'h4CE1; w_imag[873] = 16'h6657;
w_real[874] = 16'h4D81; w_imag[874] = 16'h65DD;
w_real[875] = 16'h4E21; w_imag[875] = 16'h6563;
w_real[876] = 16'h4EBF; w_imag[876] = 16'h64E8;
w_real[877] = 16'h4F5E; w_imag[877] = 16'h646C;
w_real[878] = 16'h4FFB; w_imag[878] = 16'h63EF;
w_real[879] = 16'h5097; w_imag[879] = 16'h6371;
w_real[880] = 16'h5133; w_imag[880] = 16'h62F2;
w_real[881] = 16'h51CE; w_imag[881] = 16'h6271;
w_real[882] = 16'h5269; w_imag[882] = 16'h61F1;
w_real[883] = 16'h5302; w_imag[883] = 16'h616F;
w_real[884] = 16'h539B; w_imag[884] = 16'h60EC;
w_real[885] = 16'h5433; w_imag[885] = 16'h6068;
w_real[886] = 16'h54CA; w_imag[886] = 16'h5FE3;
w_real[887] = 16'h5560; w_imag[887] = 16'h5F5E;
w_real[888] = 16'h55F5; w_imag[888] = 16'h5ED7;
w_real[889] = 16'h568A; w_imag[889] = 16'h5E50;
w_real[890] = 16'h571D; w_imag[890] = 16'h5DC7;
w_real[891] = 16'h57B0; w_imag[891] = 16'h5D3E;
w_real[892] = 16'h5842; w_imag[892] = 16'h5CB4;
w_real[893] = 16'h58D4; w_imag[893] = 16'h5C29;
w_real[894] = 16'h5964; w_imag[894] = 16'h5B9D;
w_real[895] = 16'h59F3; w_imag[895] = 16'h5B10;
w_real[896] = 16'h5A82; w_imag[896] = 16'h5A82;
w_real[897] = 16'h5B10; w_imag[897] = 16'h59F3;
w_real[898] = 16'h5B9D; w_imag[898] = 16'h5964;
w_real[899] = 16'h5C29; w_imag[899] = 16'h58D4;
w_real[900] = 16'h5CB4; w_imag[900] = 16'h5842;
w_real[901] = 16'h5D3E; w_imag[901] = 16'h57B0;
w_real[902] = 16'h5DC7; w_imag[902] = 16'h571D;
w_real[903] = 16'h5E50; w_imag[903] = 16'h568A;
w_real[904] = 16'h5ED7; w_imag[904] = 16'h55F5;
w_real[905] = 16'h5F5E; w_imag[905] = 16'h5560;
w_real[906] = 16'h5FE3; w_imag[906] = 16'h54CA;
w_real[907] = 16'h6068; w_imag[907] = 16'h5433;
w_real[908] = 16'h60EC; w_imag[908] = 16'h539B;
w_real[909] = 16'h616F; w_imag[909] = 16'h5302;
w_real[910] = 16'h61F1; w_imag[910] = 16'h5269;
w_real[911] = 16'h6271; w_imag[911] = 16'h51CE;
w_real[912] = 16'h62F2; w_imag[912] = 16'h5133;
w_real[913] = 16'h6371; w_imag[913] = 16'h5097;
w_real[914] = 16'h63EF; w_imag[914] = 16'h4FFB;
w_real[915] = 16'h646C; w_imag[915] = 16'h4F5E;
w_real[916] = 16'h64E8; w_imag[916] = 16'h4EBF;
w_real[917] = 16'h6563; w_imag[917] = 16'h4E21;
w_real[918] = 16'h65DD; w_imag[918] = 16'h4D81;
w_real[919] = 16'h6657; w_imag[919] = 16'h4CE1;
w_real[920] = 16'h66CF; w_imag[920] = 16'h4C3F;
w_real[921] = 16'h6746; w_imag[921] = 16'h4B9E;
w_real[922] = 16'h67BD; w_imag[922] = 16'h4AFB;
w_real[923] = 16'h6832; w_imag[923] = 16'h4A58;
w_real[924] = 16'h68A6; w_imag[924] = 16'h49B4;
w_real[925] = 16'h6919; w_imag[925] = 16'h490F;
w_real[926] = 16'h698C; w_imag[926] = 16'h4869;
w_real[927] = 16'h69FD; w_imag[927] = 16'h47C3;
w_real[928] = 16'h6A6D; w_imag[928] = 16'h471C;
w_real[929] = 16'h6ADC; w_imag[929] = 16'h4675;
w_real[930] = 16'h6B4A; w_imag[930] = 16'h45CD;
w_real[931] = 16'h6BB8; w_imag[931] = 16'h4524;
w_real[932] = 16'h6C24; w_imag[932] = 16'h447A;
w_real[933] = 16'h6C8F; w_imag[933] = 16'h43D0;
w_real[934] = 16'h6CF9; w_imag[934] = 16'h4325;
w_real[935] = 16'h6D62; w_imag[935] = 16'h427A;
w_real[936] = 16'h6DCA; w_imag[936] = 16'h41CE;
w_real[937] = 16'h6E30; w_imag[937] = 16'h4121;
w_real[938] = 16'h6E96; w_imag[938] = 16'h4073;
w_real[939] = 16'h6EFB; w_imag[939] = 16'h3FC5;
w_real[940] = 16'h6F5F; w_imag[940] = 16'h3F17;
w_real[941] = 16'h6FC1; w_imag[941] = 16'h3E68;
w_real[942] = 16'h7023; w_imag[942] = 16'h3DB8;
w_real[943] = 16'h7083; w_imag[943] = 16'h3D07;
w_real[944] = 16'h70E2; w_imag[944] = 16'h3C56;
w_real[945] = 16'h7141; w_imag[945] = 16'h3BA5;
w_real[946] = 16'h719E; w_imag[946] = 16'h3AF2;
w_real[947] = 16'h71FA; w_imag[947] = 16'h3A40;
w_real[948] = 16'h7255; w_imag[948] = 16'h398C;
w_real[949] = 16'h72AF; w_imag[949] = 16'h38D8;
w_real[950] = 16'h7307; w_imag[950] = 16'h3824;
w_real[951] = 16'h735F; w_imag[951] = 16'h376F;
w_real[952] = 16'h73B5; w_imag[952] = 16'h36BA;
w_real[953] = 16'h740B; w_imag[953] = 16'h3604;
w_real[954] = 16'h745F; w_imag[954] = 16'h354D;
w_real[955] = 16'h74B2; w_imag[955] = 16'h3496;
w_real[956] = 16'h7504; w_imag[956] = 16'h33DE;
w_real[957] = 16'h7555; w_imag[957] = 16'h3326;
w_real[958] = 16'h75A5; w_imag[958] = 16'h326E;
w_real[959] = 16'h75F4; w_imag[959] = 16'h31B5;
w_real[960] = 16'h7641; w_imag[960] = 16'h30FB;
w_real[961] = 16'h768E; w_imag[961] = 16'h3041;
w_real[962] = 16'h76D9; w_imag[962] = 16'h2F87;
w_real[963] = 16'h7723; w_imag[963] = 16'h2ECC;
w_real[964] = 16'h776C; w_imag[964] = 16'h2E11;
w_real[965] = 16'h77B4; w_imag[965] = 16'h2D55;
w_real[966] = 16'h77FA; w_imag[966] = 16'h2C98;
w_real[967] = 16'h7840; w_imag[967] = 16'h2BDC;
w_real[968] = 16'h7884; w_imag[968] = 16'h2B1F;
w_real[969] = 16'h78C7; w_imag[969] = 16'h2A61;
w_real[970] = 16'h7909; w_imag[970] = 16'h29A3;
w_real[971] = 16'h794A; w_imag[971] = 16'h28E5;
w_real[972] = 16'h798A; w_imag[972] = 16'h2826;
w_real[973] = 16'h79C8; w_imag[973] = 16'h2767;
w_real[974] = 16'h7A05; w_imag[974] = 16'h26A8;
w_real[975] = 16'h7A42; w_imag[975] = 16'h25E8;
w_real[976] = 16'h7A7D; w_imag[976] = 16'h2528;
w_real[977] = 16'h7AB6; w_imag[977] = 16'h2467;
w_real[978] = 16'h7AEF; w_imag[978] = 16'h23A6;
w_real[979] = 16'h7B26; w_imag[979] = 16'h22E5;
w_real[980] = 16'h7B5D; w_imag[980] = 16'h2223;
w_real[981] = 16'h7B92; w_imag[981] = 16'h2161;
w_real[982] = 16'h7BC5; w_imag[982] = 16'h209F;
w_real[983] = 16'h7BF8; w_imag[983] = 16'h1FDC;
w_real[984] = 16'h7C29; w_imag[984] = 16'h1F19;
w_real[985] = 16'h7C5A; w_imag[985] = 16'h1E56;
w_real[986] = 16'h7C89; w_imag[986] = 16'h1D93;
w_real[987] = 16'h7CB7; w_imag[987] = 16'h1CCF;
w_real[988] = 16'h7CE3; w_imag[988] = 16'h1C0B;
w_real[989] = 16'h7D0F; w_imag[989] = 16'h1B47;
w_real[990] = 16'h7D39; w_imag[990] = 16'h1A82;
w_real[991] = 16'h7D62; w_imag[991] = 16'h19BD;
w_real[992] = 16'h7D8A; w_imag[992] = 16'h18F8;
w_real[993] = 16'h7DB0; w_imag[993] = 16'h1833;
w_real[994] = 16'h7DD6; w_imag[994] = 16'h176D;
w_real[995] = 16'h7DFA; w_imag[995] = 16'h16A8;
w_real[996] = 16'h7E1D; w_imag[996] = 16'h15E2;
w_real[997] = 16'h7E3F; w_imag[997] = 16'h151B;
w_real[998] = 16'h7E5F; w_imag[998] = 16'h1455;
w_real[999] = 16'h7E7F; w_imag[999] = 16'h138E;
w_real[1000] = 16'h7E9D; w_imag[1000] = 16'h12C8;
w_real[1001] = 16'h7EBA; w_imag[1001] = 16'h1201;
w_real[1002] = 16'h7ED5; w_imag[1002] = 16'h1139;
w_real[1003] = 16'h7EF0; w_imag[1003] = 16'h1072;
w_real[1004] = 16'h7F09; w_imag[1004] = 16'h0FAB;
w_real[1005] = 16'h7F21; w_imag[1005] = 16'h0EE3;
w_real[1006] = 16'h7F38; w_imag[1006] = 16'h0E1B;
w_real[1007] = 16'h7F4D; w_imag[1007] = 16'h0D53;
w_real[1008] = 16'h7F62; w_imag[1008] = 16'h0C8B;
w_real[1009] = 16'h7F75; w_imag[1009] = 16'h0BC3;
w_real[1010] = 16'h7F87; w_imag[1010] = 16'h0AFB;
w_real[1011] = 16'h7F97; w_imag[1011] = 16'h0A33;
w_real[1012] = 16'h7FA7; w_imag[1012] = 16'h096A;
w_real[1013] = 16'h7FB5; w_imag[1013] = 16'h08A2;
w_real[1014] = 16'h7FC2; w_imag[1014] = 16'h07D9;
w_real[1015] = 16'h7FCE; w_imag[1015] = 16'h0710;
w_real[1016] = 16'h7FD8; w_imag[1016] = 16'h0647;
w_real[1017] = 16'h7FE1; w_imag[1017] = 16'h057F;
w_real[1018] = 16'h7FE9; w_imag[1018] = 16'h04B6;
w_real[1019] = 16'h7FF0; w_imag[1019] = 16'h03ED;
w_real[1020] = 16'h7FF6; w_imag[1020] = 16'h0324;
w_real[1021] = 16'h7FFA; w_imag[1021] = 16'h025B;
w_real[1022] = 16'h7FFD; w_imag[1022] = 16'h0192;
w_real[1023] = 16'h7FFF; w_imag[1023] = 16'h00C9;
