w_real[0] = 12'h7FF; w_imag[0] = 12'h000;
w_real[1] = 12'h7F6; w_imag[1] = 12'hF38;
w_real[2] = 12'h7D8; w_imag[2] = 12'hE71;
w_real[3] = 12'h7A7; w_imag[3] = 12'hDAE;
w_real[4] = 12'h764; w_imag[4] = 12'hCF1;
w_real[5] = 12'h70E; w_imag[5] = 12'hC3B;
w_real[6] = 12'h6A6; w_imag[6] = 12'hB8F;
w_real[7] = 12'h62F; w_imag[7] = 12'hAED;
w_real[8] = 12'h5A8; w_imag[8] = 12'hA58;
w_real[9] = 12'h513; w_imag[9] = 12'h9D1;
w_real[10] = 12'h471; w_imag[10] = 12'h95A;
w_real[11] = 12'h3C5; w_imag[11] = 12'h8F2;
w_real[12] = 12'h30F; w_imag[12] = 12'h89C;
w_real[13] = 12'h252; w_imag[13] = 12'h859;
w_real[14] = 12'h18F; w_imag[14] = 12'h828;
w_real[15] = 12'h0C8; w_imag[15] = 12'h80A;
w_real[16] = 12'h000; w_imag[16] = 12'h800;
w_real[17] = 12'hF38; w_imag[17] = 12'h80A;
w_real[18] = 12'hE71; w_imag[18] = 12'h828;
w_real[19] = 12'hDAE; w_imag[19] = 12'h859;
w_real[20] = 12'hCF1; w_imag[20] = 12'h89C;
w_real[21] = 12'hC3B; w_imag[21] = 12'h8F2;
w_real[22] = 12'hB8F; w_imag[22] = 12'h95A;
w_real[23] = 12'hAED; w_imag[23] = 12'h9D1;
w_real[24] = 12'hA58; w_imag[24] = 12'hA58;
w_real[25] = 12'h9D1; w_imag[25] = 12'hAED;
w_real[26] = 12'h95A; w_imag[26] = 12'hB8F;
w_real[27] = 12'h8F2; w_imag[27] = 12'hC3B;
w_real[28] = 12'h89C; w_imag[28] = 12'hCF1;
w_real[29] = 12'h859; w_imag[29] = 12'hDAE;
w_real[30] = 12'h828; w_imag[30] = 12'hE71;
w_real[31] = 12'h80A; w_imag[31] = 12'hF38;
w_real[32] = 12'h800; w_imag[32] = 12'h000;
w_real[33] = 12'h80A; w_imag[33] = 12'h0C8;
w_real[34] = 12'h828; w_imag[34] = 12'h18F;
w_real[35] = 12'h859; w_imag[35] = 12'h252;
w_real[36] = 12'h89C; w_imag[36] = 12'h30F;
w_real[37] = 12'h8F2; w_imag[37] = 12'h3C5;
w_real[38] = 12'h95A; w_imag[38] = 12'h471;
w_real[39] = 12'h9D1; w_imag[39] = 12'h513;
w_real[40] = 12'hA58; w_imag[40] = 12'h5A8;
w_real[41] = 12'hAED; w_imag[41] = 12'h62F;
w_real[42] = 12'hB8F; w_imag[42] = 12'h6A6;
w_real[43] = 12'hC3B; w_imag[43] = 12'h70E;
w_real[44] = 12'hCF1; w_imag[44] = 12'h764;
w_real[45] = 12'hDAE; w_imag[45] = 12'h7A7;
w_real[46] = 12'hE71; w_imag[46] = 12'h7D8;
w_real[47] = 12'hF38; w_imag[47] = 12'h7F6;
w_real[48] = 12'h000; w_imag[48] = 12'h7FF;
w_real[49] = 12'h0C8; w_imag[49] = 12'h7F6;
w_real[50] = 12'h18F; w_imag[50] = 12'h7D8;
w_real[51] = 12'h252; w_imag[51] = 12'h7A7;
w_real[52] = 12'h30F; w_imag[52] = 12'h764;
w_real[53] = 12'h3C5; w_imag[53] = 12'h70E;
w_real[54] = 12'h471; w_imag[54] = 12'h6A6;
w_real[55] = 12'h513; w_imag[55] = 12'h62F;
w_real[56] = 12'h5A8; w_imag[56] = 12'h5A8;
w_real[57] = 12'h62F; w_imag[57] = 12'h513;
w_real[58] = 12'h6A6; w_imag[58] = 12'h471;
w_real[59] = 12'h70E; w_imag[59] = 12'h3C5;
w_real[60] = 12'h764; w_imag[60] = 12'h30F;
w_real[61] = 12'h7A7; w_imag[61] = 12'h252;
w_real[62] = 12'h7D8; w_imag[62] = 12'h18F;
w_real[63] = 12'h7F6; w_imag[63] = 12'h0C8;
