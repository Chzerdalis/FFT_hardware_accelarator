0 0
77 -1584
320 -3253
821 -5536
1594 -8014
3233 -12909
3009 -9920
4506 -12594
6469 -15618
9211 -19476
13361 -24998
21172 -35324
75161 -112486
11937 -16095
36224 -44139
125355 -138308
130035 -130035
152429 -138153
50467 -41417
-51918 38505
-49736 33233
-73406 43997
-22680 12123
-71072 33614
-47509 19679
-53211 19039
-44499 13498
-44479 11141
-42454 8444
-42871 6359
-41083 4046
-40379 1983
-40174 0
-40379 -1983
-41083 -4046
-42871 -6359
-42454 -8444
-44479 -11141
-44499 -13498
-53211 -19039
-47509 -19679
-71072 -33614
-22680 -12123
-73406 -43997
-49736 -33233
-51918 -38505
50467 41417
152429 138153
130035 130035
125355 138308
36224 44139
11937 16095
75161 112486
21172 35324
13361 24998
9211 19476
6469 15618
4506 12594
3009 9920
3233 12909
1594 8014
821 5536
320 3253
77 1584
