gen_input_real[0] = 18'sd0;
gen_input_real[256] = 18'sd255;
gen_input_real[512] = -18'sd16;
gen_input_real[768] = -18'sd150;
gen_input_real[64] = 18'sd7;
gen_input_real[320] = 18'sd67;
gen_input_real[576] = 18'sd19;
gen_input_real[832] = -18'sd54;
gen_input_real[128] = -18'sd32;
gen_input_real[384] = 18'sd70;
gen_input_real[640] = 18'sd16;
gen_input_real[896] = -18'sd83;
gen_input_real[192] = 18'sd15;
gen_input_real[448] = 18'sd82;
gen_input_real[704] = -18'sd33;
gen_input_real[960] = -18'sd60;
gen_input_real[16] = 18'sd18;
gen_input_real[272] = 18'sd40;
gen_input_real[528] = 18'sd9;
gen_input_real[784] = -18'sd52;
gen_input_real[80] = -18'sd22;
gen_input_real[336] = 18'sd75;
gen_input_real[592] = 18'sd11;
gen_input_real[848] = -18'sd65;
gen_input_real[144] = 18'sd16;
gen_input_real[400] = 18'sd34;
gen_input_real[656] = -18'sd31;
gen_input_real[912] = -18'sd20;
gen_input_real[208] = 18'sd6;
gen_input_real[464] = 18'sd30;
gen_input_real[720] = 18'sd36;
gen_input_real[976] = -18'sd56;
gen_input_real[32] = -18'sd67;
gen_input_real[288] = 18'sd92;
gen_input_real[544] = 18'sd87;
gen_input_real[800] = -18'sd120;
gen_input_real[96] = -18'sd103;
gen_input_real[352] = 18'sd115;
gen_input_real[608] = 18'sd107;
gen_input_real[864] = -18'sd93;
gen_input_real[160] = -18'sd101;
gen_input_real[416] = 18'sd91;
gen_input_real[672] = 18'sd90;
gen_input_real[928] = -18'sd104;
gen_input_real[224] = -18'sd77;
gen_input_real[480] = 18'sd89;
gen_input_real[736] = 18'sd70;
gen_input_real[992] = -18'sd44;
gen_input_real[48] = -18'sd76;
gen_input_real[304] = 18'sd14;
gen_input_real[560] = 18'sd72;
gen_input_real[816] = -18'sd32;
gen_input_real[112] = -18'sd39;
gen_input_real[368] = 18'sd77;
gen_input_real[624] = 18'sd2;
gen_input_real[880] = -18'sd105;
gen_input_real[176] = 18'sd4;
gen_input_real[432] = 18'sd104;
gen_input_real[688] = 18'sd12;
gen_input_real[944] = -18'sd93;
gen_input_real[240] = -18'sd17;
gen_input_real[496] = 18'sd88;
gen_input_real[752] = 18'sd11;
gen_input_real[1008] = -18'sd75;
gen_input_real[4] = -18'sd9;
gen_input_real[260] = 18'sd48;
gen_input_real[516] = 18'sd11;
gen_input_real[772] = -18'sd23;
gen_input_real[68] = -18'sd18;
gen_input_real[324] = 18'sd5;
gen_input_real[580] = 18'sd35;
gen_input_real[836] = -18'sd6;
gen_input_real[132] = -18'sd58;
gen_input_real[388] = 18'sd29;
gen_input_real[644] = 18'sd81;
gen_input_real[900] = -18'sd43;
gen_input_real[196] = -18'sd107;
gen_input_real[452] = 18'sd32;
gen_input_real[708] = 18'sd128;
gen_input_real[964] = -18'sd9;
gen_input_real[20] = -18'sd116;
gen_input_real[276] = -18'sd17;
gen_input_real[532] = 18'sd81;
gen_input_real[788] = 18'sd48;
gen_input_real[84] = -18'sd55;
gen_input_real[340] = -18'sd65;
gen_input_real[596] = 18'sd38;
gen_input_real[852] = 18'sd42;
gen_input_real[148] = -18'sd32;
gen_input_real[404] = 18'sd10;
gen_input_real[660] = 18'sd60;
gen_input_real[916] = -18'sd55;
gen_input_real[212] = -18'sd98;
gen_input_real[468] = 18'sd76;
gen_input_real[724] = 18'sd96;
gen_input_real[980] = -18'sd80;
gen_input_real[36] = -18'sd68;
gen_input_real[292] = 18'sd74;
gen_input_real[548] = 18'sd49;
gen_input_real[804] = -18'sd64;
gen_input_real[100] = -18'sd52;
gen_input_real[356] = 18'sd53;
gen_input_real[612] = 18'sd60;
gen_input_real[868] = -18'sd53;
gen_input_real[164] = -18'sd53;
gen_input_real[420] = 18'sd58;
gen_input_real[676] = 18'sd28;
gen_input_real[932] = -18'sd40;
gen_input_real[228] = -18'sd6;
gen_input_real[484] = 18'sd4;
gen_input_real[740] = 18'sd28;
gen_input_real[996] = 18'sd17;
gen_input_real[52] = -18'sd78;
gen_input_real[308] = -18'sd20;
gen_input_real[564] = 18'sd87;
gen_input_real[820] = 18'sd13;
gen_input_real[116] = -18'sd36;
gen_input_real[372] = -18'sd8;
gen_input_real[628] = -18'sd17;
gen_input_real[884] = 18'sd19;
gen_input_real[180] = 18'sd34;
gen_input_real[436] = -18'sd47;
gen_input_real[692] = -18'sd21;
gen_input_real[948] = 18'sd70;
gen_input_real[244] = 18'sd6;
gen_input_real[500] = -18'sd67;
gen_input_real[756] = 18'sd8;
gen_input_real[1012] = 18'sd46;
gen_input_real[8] = -18'sd21;
gen_input_real[264] = -18'sd23;
gen_input_real[520] = 18'sd29;
gen_input_real[776] = 18'sd0;
gen_input_real[72] = -18'sd42;
gen_input_real[328] = 18'sd24;
gen_input_real[584] = 18'sd72;
gen_input_real[840] = -18'sd35;
gen_input_real[136] = -18'sd102;
gen_input_real[392] = 18'sd21;
gen_input_real[648] = 18'sd109;
gen_input_real[904] = 18'sd3;
gen_input_real[200] = -18'sd90;
gen_input_real[456] = -18'sd18;
gen_input_real[712] = 18'sd58;
gen_input_real[968] = 18'sd19;
gen_input_real[24] = -18'sd29;
gen_input_real[280] = -18'sd12;
gen_input_real[536] = 18'sd20;
gen_input_real[792] = 18'sd2;
gen_input_real[88] = -18'sd30;
gen_input_real[344] = 18'sd2;
gen_input_real[600] = 18'sd36;
gen_input_real[856] = -18'sd5;
gen_input_real[152] = -18'sd32;
gen_input_real[408] = 18'sd15;
gen_input_real[664] = 18'sd24;
gen_input_real[920] = -18'sd29;
gen_input_real[216] = -18'sd10;
gen_input_real[472] = 18'sd34;
gen_input_real[728] = -18'sd26;
gen_input_real[984] = -18'sd19;
gen_input_real[40] = 18'sd89;
gen_input_real[296] = -18'sd5;
gen_input_real[552] = -18'sd124;
gen_input_real[808] = 18'sd12;
gen_input_real[104] = 18'sd85;
gen_input_real[360] = 18'sd12;
gen_input_real[616] = -18'sd14;
gen_input_real[872] = -18'sd46;
gen_input_real[168] = -18'sd21;
gen_input_real[424] = 18'sd41;
gen_input_real[680] = 18'sd24;
gen_input_real[936] = 18'sd0;
gen_input_real[232] = -18'sd27;
gen_input_real[488] = -18'sd36;
gen_input_real[744] = 18'sd31;
gen_input_real[1000] = 18'sd55;
gen_input_real[56] = -18'sd24;
gen_input_real[312] = -18'sd52;
gen_input_real[568] = 18'sd15;
gen_input_real[824] = 18'sd28;
gen_input_real[120] = -18'sd3;
gen_input_real[376] = -18'sd16;
gen_input_real[632] = -18'sd15;
gen_input_real[888] = 18'sd34;
gen_input_real[184] = 18'sd14;
gen_input_real[440] = -18'sd52;
gen_input_real[696] = 18'sd11;
gen_input_real[952] = 18'sd41;
gen_input_real[248] = -18'sd29;
gen_input_real[504] = -18'sd8;
gen_input_real[760] = 18'sd33;
gen_input_real[1016] = -18'sd27;
gen_input_real[12] = -18'sd29;
gen_input_real[268] = 18'sd55;
gen_input_real[524] = 18'sd14;
gen_input_real[780] = -18'sd70;
gen_input_real[76] = 18'sd11;
gen_input_real[332] = 18'sd72;
gen_input_real[588] = -18'sd29;
gen_input_real[844] = -18'sd78;
gen_input_real[140] = 18'sd19;
gen_input_real[396] = 18'sd90;
gen_input_real[652] = 18'sd0;
gen_input_real[908] = -18'sd83;
gen_input_real[204] = 18'sd4;
gen_input_real[460] = 18'sd55;
gen_input_real[716] = -18'sd15;
gen_input_real[972] = -18'sd33;
gen_input_real[28] = -18'sd1;
gen_input_real[284] = 18'sd43;
gen_input_real[540] = 18'sd29;
gen_input_real[796] = -18'sd64;
gen_input_real[92] = -18'sd30;
gen_input_real[348] = 18'sd50;
gen_input_real[604] = -18'sd4;
gen_input_real[860] = -18'sd4;
gen_input_real[156] = 18'sd46;
gen_input_real[412] = -18'sd28;
gen_input_real[668] = -18'sd73;
gen_input_real[924] = 18'sd25;
gen_input_real[220] = 18'sd82;
gen_input_real[476] = -18'sd1;
gen_input_real[732] = -18'sd73;
gen_input_real[988] = -18'sd24;
gen_input_real[44] = 18'sd53;
gen_input_real[300] = 18'sd39;
gen_input_real[556] = -18'sd26;
gen_input_real[812] = -18'sd33;
gen_input_real[108] = -18'sd5;
gen_input_real[364] = 18'sd15;
gen_input_real[620] = 18'sd39;
gen_input_real[876] = -18'sd12;
gen_input_real[172] = -18'sd63;
gen_input_real[428] = 18'sd34;
gen_input_real[684] = 18'sd59;
gen_input_real[940] = -18'sd65;
gen_input_real[236] = -18'sd33;
gen_input_real[492] = 18'sd82;
gen_input_real[748] = 18'sd10;
gen_input_real[1004] = -18'sd81;
gen_input_real[60] = -18'sd11;
gen_input_real[316] = 18'sd64;
gen_input_real[572] = 18'sd37;
gen_input_real[828] = -18'sd39;
gen_input_real[124] = -18'sd82;
gen_input_real[380] = 18'sd39;
gen_input_real[636] = 18'sd123;
gen_input_real[892] = -18'sd66;
gen_input_real[188] = -18'sd113;
gen_input_real[444] = 18'sd68;
gen_input_real[700] = 18'sd42;
gen_input_real[956] = -18'sd39;
gen_input_real[252] = 18'sd26;
gen_input_real[508] = 18'sd40;
gen_input_real[764] = -18'sd42;
gen_input_real[1020] = -18'sd80;
gen_input_real[1] = 18'sd25;
gen_input_real[257] = 18'sd113;
gen_input_real[513] = -18'sd12;
gen_input_real[769] = -18'sd118;
gen_input_real[65] = 18'sd18;
gen_input_real[321] = 18'sd111;
gen_input_real[577] = -18'sd32;
gen_input_real[833] = -18'sd88;
gen_input_real[129] = 18'sd29;
gen_input_real[385] = 18'sd53;
gen_input_real[641] = 18'sd0;
gen_input_real[897] = -18'sd39;
gen_input_real[193] = -18'sd47;
gen_input_real[449] = 18'sd49;
gen_input_real[705] = 18'sd80;
gen_input_real[961] = -18'sd60;
gen_input_real[17] = -18'sd70;
gen_input_real[273] = 18'sd67;
gen_input_real[529] = 18'sd35;
gen_input_real[785] = -18'sd58;
gen_input_real[81] = -18'sd20;
gen_input_real[337] = 18'sd20;
gen_input_real[593] = 18'sd38;
gen_input_real[849] = 18'sd18;
gen_input_real[145] = -18'sd64;
gen_input_real[401] = -18'sd20;
gen_input_real[657] = 18'sd81;
gen_input_real[913] = -18'sd4;
gen_input_real[209] = -18'sd89;
gen_input_real[465] = 18'sd15;
gen_input_real[721] = 18'sd85;
gen_input_real[977] = -18'sd10;
gen_input_real[33] = -18'sd77;
gen_input_real[289] = 18'sd19;
gen_input_real[545] = 18'sd86;
gen_input_real[801] = -18'sd47;
gen_input_real[97] = -18'sd94;
gen_input_real[353] = 18'sd71;
gen_input_real[609] = 18'sd70;
gen_input_real[865] = -18'sd88;
gen_input_real[161] = -18'sd37;
gen_input_real[417] = 18'sd106;
gen_input_real[673] = 18'sd33;
gen_input_real[929] = -18'sd123;
gen_input_real[225] = -18'sd61;
gen_input_real[481] = 18'sd126;
gen_input_real[737] = 18'sd98;
gen_input_real[993] = -18'sd103;
gen_input_real[49] = -18'sd127;
gen_input_real[305] = 18'sd59;
gen_input_real[561] = 18'sd133;
gen_input_real[817] = -18'sd23;
gen_input_real[113] = -18'sd109;
gen_input_real[369] = 18'sd23;
gen_input_real[625] = 18'sd73;
gen_input_real[881] = -18'sd42;
gen_input_real[177] = -18'sd48;
gen_input_real[433] = 18'sd47;
gen_input_real[689] = 18'sd38;
gen_input_real[945] = -18'sd37;
gen_input_real[241] = -18'sd26;
gen_input_real[497] = 18'sd26;
gen_input_real[753] = 18'sd19;
gen_input_real[1009] = -18'sd9;
gen_input_real[5] = -18'sd31;
gen_input_real[261] = -18'sd21;
gen_input_real[517] = 18'sd56;
gen_input_real[773] = 18'sd47;
gen_input_real[69] = -18'sd76;
gen_input_real[325] = -18'sd52;
gen_input_real[581] = 18'sd80;
gen_input_real[837] = 18'sd30;
gen_input_real[133] = -18'sd66;
gen_input_real[389] = 18'sd5;
gen_input_real[645] = 18'sd55;
gen_input_real[901] = -18'sd31;
gen_input_real[197] = -18'sd74;
gen_input_real[453] = 18'sd40;
gen_input_real[709] = 18'sd108;
gen_input_real[965] = -18'sd40;
gen_input_real[21] = -18'sd134;
gen_input_real[277] = 18'sd26;
gen_input_real[533] = 18'sd154;
gen_input_real[789] = 18'sd3;
gen_input_real[85] = -18'sd164;
gen_input_real[341] = -18'sd27;
gen_input_real[597] = 18'sd147;
gen_input_real[853] = 18'sd33;
gen_input_real[149] = -18'sd126;
gen_input_real[405] = -18'sd24;
gen_input_real[661] = 18'sd129;
gen_input_real[917] = 18'sd14;
gen_input_real[213] = -18'sd138;
gen_input_real[469] = -18'sd12;
gen_input_real[725] = 18'sd123;
gen_input_real[981] = 18'sd1;
gen_input_real[37] = -18'sd94;
gen_input_real[293] = 18'sd27;
gen_input_real[549] = 18'sd55;
gen_input_real[805] = -18'sd47;
gen_input_real[101] = -18'sd8;
gen_input_real[357] = 18'sd30;
gen_input_real[613] = 18'sd0;
gen_input_real[869] = 18'sd8;
gen_input_real[165] = -18'sd43;
gen_input_real[421] = -18'sd32;
gen_input_real[677] = 18'sd75;
gen_input_real[933] = 18'sd19;
gen_input_real[229] = -18'sd67;
gen_input_real[485] = 18'sd5;
gen_input_real[741] = 18'sd55;
gen_input_real[997] = -18'sd8;
gen_input_real[53] = -18'sd60;
gen_input_real[309] = -18'sd19;
gen_input_real[565] = 18'sd60;
gen_input_real[821] = 18'sd45;
gen_input_real[117] = -18'sd54;
gen_input_real[373] = -18'sd44;
gen_input_real[629] = 18'sd68;
gen_input_real[885] = 18'sd39;
gen_input_real[181] = -18'sd94;
gen_input_real[437] = -18'sd52;
gen_input_real[693] = 18'sd98;
gen_input_real[949] = 18'sd81;
gen_input_real[245] = -18'sd91;
gen_input_real[501] = -18'sd123;
gen_input_real[757] = 18'sd96;
gen_input_real[1013] = 18'sd161;
gen_input_real[9] = -18'sd97;
gen_input_real[265] = -18'sd154;
gen_input_real[521] = 18'sd80;
gen_input_real[777] = 18'sd99;
gen_input_real[73] = -18'sd62;
gen_input_real[329] = -18'sd35;
gen_input_real[585] = 18'sd57;
gen_input_real[841] = -18'sd6;
gen_input_real[137] = -18'sd57;
gen_input_real[393] = 18'sd17;
gen_input_real[649] = 18'sd67;
gen_input_real[905] = -18'sd2;
gen_input_real[201] = -18'sd83;
gen_input_real[457] = -18'sd25;
gen_input_real[713] = 18'sd82;
gen_input_real[969] = 18'sd42;
gen_input_real[25] = -18'sd64;
gen_input_real[281] = -18'sd39;
gen_input_real[537] = 18'sd63;
gen_input_real[793] = 18'sd32;
gen_input_real[89] = -18'sd81;
gen_input_real[345] = -18'sd24;
gen_input_real[601] = 18'sd80;
gen_input_real[857] = 18'sd1;
gen_input_real[153] = -18'sd45;
gen_input_real[409] = 18'sd13;
gen_input_real[665] = 18'sd19;
gen_input_real[921] = 18'sd16;
gen_input_real[217] = -18'sd32;
gen_input_real[473] = -18'sd65;
gen_input_real[729] = 18'sd53;
gen_input_real[985] = 18'sd89;
gen_input_real[41] = -18'sd31;
gen_input_real[297] = -18'sd95;
gen_input_real[553] = -18'sd26;
gen_input_real[809] = 18'sd106;
gen_input_real[105] = 18'sd62;
gen_input_real[361] = -18'sd112;
gen_input_real[617] = -18'sd53;
gen_input_real[873] = 18'sd107;
gen_input_real[169] = 18'sd17;
gen_input_real[425] = -18'sd100;
gen_input_real[681] = 18'sd24;
gen_input_real[937] = 18'sd75;
gen_input_real[233] = -18'sd41;
gen_input_real[489] = -18'sd31;
gen_input_real[745] = 18'sd20;
gen_input_real[1001] = 18'sd14;
gen_input_real[57] = 18'sd3;
gen_input_real[313] = -18'sd40;
gen_input_real[569] = 18'sd8;
gen_input_real[825] = 18'sd70;
gen_input_real[121] = -18'sd48;
gen_input_real[377] = -18'sd80;
gen_input_real[633] = 18'sd84;
gen_input_real[889] = 18'sd81;
gen_input_real[185] = -18'sd95;
gen_input_real[441] = -18'sd75;
gen_input_real[697] = 18'sd77;
gen_input_real[953] = 18'sd68;
gen_input_real[249] = -18'sd47;
gen_input_real[505] = -18'sd67;
gen_input_real[761] = 18'sd33;
gen_input_real[1017] = 18'sd55;
gen_input_real[13] = -18'sd46;
gen_input_real[269] = -18'sd25;
gen_input_real[525] = 18'sd49;
gen_input_real[781] = -18'sd2;
gen_input_real[77] = -18'sd10;
gen_input_real[333] = 18'sd1;
gen_input_real[589] = -18'sd41;
gen_input_real[845] = 18'sd24;
gen_input_real[141] = 18'sd53;
gen_input_real[397] = -18'sd49;
gen_input_real[653] = -18'sd25;
gen_input_real[909] = 18'sd51;
gen_input_real[205] = 18'sd20;
gen_input_real[461] = -18'sd31;
gen_input_real[717] = -18'sd59;
gen_input_real[973] = 18'sd5;
gen_input_real[29] = 18'sd84;
gen_input_real[285] = 18'sd13;
gen_input_real[541] = -18'sd56;
gen_input_real[797] = -18'sd21;
gen_input_real[93] = 18'sd1;
gen_input_real[349] = 18'sd20;
gen_input_real[605] = 18'sd34;
gen_input_real[861] = -18'sd2;
gen_input_real[157] = -18'sd29;
gen_input_real[413] = -18'sd36;
gen_input_real[669] = -18'sd9;
gen_input_real[925] = 18'sd84;
gen_input_real[221] = 18'sd44;
gen_input_real[477] = -18'sd120;
gen_input_real[733] = -18'sd39;
gen_input_real[989] = 18'sd130;
gen_input_real[45] = 18'sd3;
gen_input_real[301] = -18'sd105;
gen_input_real[557] = 18'sd24;
gen_input_real[813] = 18'sd58;
gen_input_real[109] = -18'sd23;
gen_input_real[365] = -18'sd19;
gen_input_real[621] = 18'sd12;
gen_input_real[877] = 18'sd17;
gen_input_real[173] = -18'sd5;
gen_input_real[429] = -18'sd37;
gen_input_real[685] = 18'sd1;
gen_input_real[941] = 18'sd42;
gen_input_real[237] = -18'sd5;
gen_input_real[493] = -18'sd20;
gen_input_real[749] = 18'sd13;
gen_input_real[1005] = -18'sd10;
gen_input_real[61] = 18'sd0;
gen_input_real[317] = 18'sd33;
gen_input_real[573] = -18'sd28;
gen_input_real[829] = -18'sd37;
gen_input_real[125] = 18'sd20;
gen_input_real[381] = 18'sd35;
gen_input_real[637] = 18'sd32;
gen_input_real[893] = -18'sd40;
gen_input_real[189] = -18'sd74;
gen_input_real[445] = 18'sd43;
gen_input_real[701] = 18'sd67;
gen_input_real[957] = -18'sd40;
gen_input_real[253] = -18'sd30;
gen_input_real[509] = 18'sd39;
gen_input_real[765] = -18'sd7;
gen_input_real[1021] = -18'sd32;
gen_input_real[2] = 18'sd32;
gen_input_real[258] = 18'sd7;
gen_input_real[514] = -18'sd39;
gen_input_real[770] = 18'sd30;
gen_input_real[66] = 18'sd40;
gen_input_real[322] = -18'sd67;
gen_input_real[578] = -18'sd43;
gen_input_real[834] = 18'sd74;
gen_input_real[130] = 18'sd40;
gen_input_real[386] = -18'sd32;
gen_input_real[642] = -18'sd35;
gen_input_real[898] = -18'sd20;
gen_input_real[194] = 18'sd37;
gen_input_real[450] = 18'sd28;
gen_input_real[706] = -18'sd33;
gen_input_real[962] = 18'sd0;
gen_input_real[18] = 18'sd10;
gen_input_real[274] = -18'sd13;
gen_input_real[530] = 18'sd20;
gen_input_real[786] = 18'sd5;
gen_input_real[82] = -18'sd42;
gen_input_real[338] = -18'sd1;
gen_input_real[594] = 18'sd37;
gen_input_real[850] = 18'sd5;
gen_input_real[146] = -18'sd17;
gen_input_real[402] = -18'sd12;
gen_input_real[658] = 18'sd19;
gen_input_real[914] = 18'sd23;
gen_input_real[210] = -18'sd58;
gen_input_real[466] = -18'sd24;
gen_input_real[722] = 18'sd105;
gen_input_real[978] = -18'sd3;
gen_input_real[34] = -18'sd130;
gen_input_real[290] = 18'sd39;
gen_input_real[546] = 18'sd120;
gen_input_real[802] = -18'sd44;
gen_input_real[98] = -18'sd84;
gen_input_real[354] = 18'sd9;
gen_input_real[610] = 18'sd36;
gen_input_real[866] = 18'sd29;
gen_input_real[162] = 18'sd2;
gen_input_real[418] = -18'sd34;
gen_input_real[674] = -18'sd20;
gen_input_real[930] = -18'sd1;
gen_input_real[226] = 18'sd21;
gen_input_real[482] = 18'sd56;
gen_input_real[738] = -18'sd13;
gen_input_real[994] = -18'sd84;
gen_input_real[50] = -18'sd5;
gen_input_real[306] = 18'sd59;
gen_input_real[562] = 18'sd31;
gen_input_real[818] = -18'sd20;
gen_input_real[114] = -18'sd51;
gen_input_real[370] = 18'sd25;
gen_input_real[626] = 18'sd49;
gen_input_real[882] = -18'sd53;
gen_input_real[178] = -18'sd24;
gen_input_real[434] = 18'sd41;
gen_input_real[690] = -18'sd1;
gen_input_real[946] = 18'sd10;
gen_input_real[242] = 18'sd2;
gen_input_real[498] = -18'sd49;
gen_input_real[754] = 18'sd25;
gen_input_real[1010] = 18'sd46;
gen_input_real[6] = -18'sd55;
gen_input_real[262] = -18'sd33;
gen_input_real[518] = 18'sd67;
gen_input_real[774] = 18'sd47;
gen_input_real[70] = -18'sd68;
gen_input_real[326] = -18'sd77;
gen_input_real[582] = 18'sd75;
gen_input_real[838] = 18'sd95;
gen_input_real[134] = -18'sd81;
gen_input_real[390] = -18'sd84;
gen_input_real[646] = 18'sd80;
gen_input_real[902] = 18'sd48;
gen_input_real[198] = -18'sd70;
gen_input_real[454] = -18'sd8;
gen_input_real[710] = 18'sd40;
gen_input_real[966] = -18'sd3;
gen_input_real[22] = -18'sd14;
gen_input_real[278] = -18'sd20;
gen_input_real[534] = 18'sd31;
gen_input_real[790] = 18'sd41;
gen_input_real[86] = -18'sd75;
gen_input_real[342] = -18'sd24;
gen_input_real[598] = 18'sd100;
gen_input_real[854] = -18'sd17;
gen_input_real[150] = -18'sd107;
gen_input_real[406] = 18'sd53;
gen_input_real[662] = 18'sd112;
gen_input_real[918] = -18'sd62;
gen_input_real[214] = -18'sd106;
gen_input_real[470] = 18'sd26;
gen_input_real[726] = 18'sd95;
gen_input_real[982] = 18'sd31;
gen_input_real[38] = -18'sd89;
gen_input_real[294] = -18'sd53;
gen_input_real[550] = 18'sd65;
gen_input_real[806] = 18'sd32;
gen_input_real[102] = -18'sd16;
gen_input_real[358] = -18'sd19;
gen_input_real[614] = -18'sd13;
gen_input_real[870] = 18'sd45;
gen_input_real[166] = -18'sd1;
gen_input_real[422] = -18'sd80;
gen_input_real[678] = 18'sd24;
gen_input_real[934] = 18'sd81;
gen_input_real[230] = -18'sd32;
gen_input_real[486] = -18'sd63;
gen_input_real[742] = 18'sd39;
gen_input_real[998] = 18'sd64;
gen_input_real[54] = -18'sd42;
gen_input_real[310] = -18'sd82;
gen_input_real[566] = 18'sd25;
gen_input_real[822] = 18'sd83;
gen_input_real[118] = 18'sd2;
gen_input_real[374] = -18'sd67;
gen_input_real[630] = -18'sd17;
gen_input_real[886] = 18'sd57;
gen_input_real[182] = 18'sd6;
gen_input_real[438] = -18'sd57;
gen_input_real[694] = 18'sd35;
gen_input_real[950] = 18'sd62;
gen_input_real[246] = -18'sd99;
gen_input_real[502] = -18'sd80;
gen_input_real[758] = 18'sd154;
gen_input_real[1014] = 18'sd97;
gen_input_real[10] = -18'sd161;
gen_input_real[266] = -18'sd96;
gen_input_real[522] = 18'sd123;
gen_input_real[778] = 18'sd91;
gen_input_real[74] = -18'sd81;
gen_input_real[330] = -18'sd98;
gen_input_real[586] = 18'sd52;
gen_input_real[842] = 18'sd94;
gen_input_real[138] = -18'sd39;
gen_input_real[394] = -18'sd68;
gen_input_real[650] = 18'sd44;
gen_input_real[906] = 18'sd54;
gen_input_real[202] = -18'sd45;
gen_input_real[458] = -18'sd60;
gen_input_real[714] = 18'sd19;
gen_input_real[970] = 18'sd60;
gen_input_real[26] = 18'sd8;
gen_input_real[282] = -18'sd55;
gen_input_real[538] = -18'sd5;
gen_input_real[794] = 18'sd67;
gen_input_real[90] = -18'sd19;
gen_input_real[346] = -18'sd75;
gen_input_real[602] = 18'sd32;
gen_input_real[858] = 18'sd43;
gen_input_real[154] = -18'sd8;
gen_input_real[410] = 18'sd0;
gen_input_real[666] = -18'sd30;
gen_input_real[922] = 18'sd8;
gen_input_real[218] = 18'sd47;
gen_input_real[474] = -18'sd55;
gen_input_real[730] = -18'sd27;
gen_input_real[986] = 18'sd94;
gen_input_real[42] = -18'sd1;
gen_input_real[298] = -18'sd123;
gen_input_real[554] = 18'sd12;
gen_input_real[810] = 18'sd138;
gen_input_real[106] = -18'sd14;
gen_input_real[362] = -18'sd129;
gen_input_real[618] = 18'sd24;
gen_input_real[874] = 18'sd126;
gen_input_real[170] = -18'sd33;
gen_input_real[426] = -18'sd147;
gen_input_real[682] = 18'sd27;
gen_input_real[938] = 18'sd164;
gen_input_real[234] = -18'sd3;
gen_input_real[490] = -18'sd154;
gen_input_real[746] = -18'sd26;
gen_input_real[1002] = 18'sd134;
gen_input_real[58] = 18'sd40;
gen_input_real[314] = -18'sd108;
gen_input_real[570] = -18'sd40;
gen_input_real[826] = 18'sd74;
gen_input_real[122] = 18'sd31;
gen_input_real[378] = -18'sd55;
gen_input_real[634] = -18'sd5;
gen_input_real[890] = 18'sd66;
gen_input_real[186] = -18'sd30;
gen_input_real[442] = -18'sd80;
gen_input_real[698] = 18'sd52;
gen_input_real[954] = 18'sd76;
gen_input_real[250] = -18'sd47;
gen_input_real[506] = -18'sd56;
gen_input_real[762] = 18'sd21;
gen_input_real[1018] = 18'sd31;
gen_input_real[14] = 18'sd9;
gen_input_real[270] = -18'sd19;
gen_input_real[526] = -18'sd26;
gen_input_real[782] = 18'sd26;
gen_input_real[78] = 18'sd37;
gen_input_real[334] = -18'sd38;
gen_input_real[590] = -18'sd47;
gen_input_real[846] = 18'sd48;
gen_input_real[142] = 18'sd42;
gen_input_real[398] = -18'sd73;
gen_input_real[654] = -18'sd23;
gen_input_real[910] = 18'sd109;
gen_input_real[206] = 18'sd23;
gen_input_real[462] = -18'sd133;
gen_input_real[718] = -18'sd59;
gen_input_real[974] = 18'sd127;
gen_input_real[30] = 18'sd103;
gen_input_real[286] = -18'sd98;
gen_input_real[542] = -18'sd126;
gen_input_real[798] = 18'sd61;
gen_input_real[94] = 18'sd123;
gen_input_real[350] = -18'sd33;
gen_input_real[606] = -18'sd106;
gen_input_real[862] = 18'sd37;
gen_input_real[158] = 18'sd88;
gen_input_real[414] = -18'sd70;
gen_input_real[670] = -18'sd71;
gen_input_real[926] = 18'sd94;
gen_input_real[222] = 18'sd47;
gen_input_real[478] = -18'sd86;
gen_input_real[734] = -18'sd19;
gen_input_real[990] = 18'sd77;
gen_input_real[46] = 18'sd10;
gen_input_real[302] = -18'sd85;
gen_input_real[558] = -18'sd15;
gen_input_real[814] = 18'sd89;
gen_input_real[110] = 18'sd4;
gen_input_real[366] = -18'sd81;
gen_input_real[622] = 18'sd20;
gen_input_real[878] = 18'sd64;
gen_input_real[174] = -18'sd18;
gen_input_real[430] = -18'sd38;
gen_input_real[686] = -18'sd20;
gen_input_real[942] = 18'sd20;
gen_input_real[238] = 18'sd58;
gen_input_real[494] = -18'sd35;
gen_input_real[750] = -18'sd67;
gen_input_real[1006] = 18'sd70;
gen_input_real[62] = 18'sd60;
gen_input_real[318] = -18'sd80;
gen_input_real[574] = -18'sd49;
gen_input_real[830] = 18'sd47;
gen_input_real[126] = 18'sd39;
gen_input_real[382] = 18'sd0;
gen_input_real[638] = -18'sd53;
gen_input_real[894] = -18'sd29;
gen_input_real[190] = 18'sd88;
gen_input_real[446] = 18'sd32;
gen_input_real[702] = -18'sd111;
gen_input_real[958] = -18'sd18;
gen_input_real[254] = 18'sd118;
gen_input_real[510] = 18'sd12;
gen_input_real[766] = -18'sd113;
gen_input_real[1022] = -18'sd25;
gen_input_real[3] = 18'sd80;
gen_input_real[259] = 18'sd42;
gen_input_real[515] = -18'sd40;
gen_input_real[771] = -18'sd26;
gen_input_real[67] = 18'sd39;
gen_input_real[323] = -18'sd42;
gen_input_real[579] = -18'sd68;
gen_input_real[835] = 18'sd113;
gen_input_real[131] = 18'sd66;
gen_input_real[387] = -18'sd123;
gen_input_real[643] = -18'sd39;
gen_input_real[899] = 18'sd82;
gen_input_real[195] = 18'sd39;
gen_input_real[451] = -18'sd37;
gen_input_real[707] = -18'sd64;
gen_input_real[963] = 18'sd11;
gen_input_real[19] = 18'sd81;
gen_input_real[275] = -18'sd10;
gen_input_real[531] = -18'sd82;
gen_input_real[787] = 18'sd33;
gen_input_real[83] = 18'sd65;
gen_input_real[339] = -18'sd59;
gen_input_real[595] = -18'sd34;
gen_input_real[851] = 18'sd63;
gen_input_real[147] = 18'sd12;
gen_input_real[403] = -18'sd39;
gen_input_real[659] = -18'sd15;
gen_input_real[915] = 18'sd5;
gen_input_real[211] = 18'sd33;
gen_input_real[467] = 18'sd26;
gen_input_real[723] = -18'sd39;
gen_input_real[979] = -18'sd53;
gen_input_real[35] = 18'sd24;
gen_input_real[291] = 18'sd73;
gen_input_real[547] = 18'sd1;
gen_input_real[803] = -18'sd82;
gen_input_real[99] = -18'sd25;
gen_input_real[355] = 18'sd73;
gen_input_real[611] = 18'sd28;
gen_input_real[867] = -18'sd46;
gen_input_real[163] = 18'sd4;
gen_input_real[419] = 18'sd4;
gen_input_real[675] = -18'sd50;
gen_input_real[931] = 18'sd30;
gen_input_real[227] = 18'sd64;
gen_input_real[483] = -18'sd29;
gen_input_real[739] = -18'sd43;
gen_input_real[995] = 18'sd1;
gen_input_real[51] = 18'sd33;
gen_input_real[307] = 18'sd15;
gen_input_real[563] = -18'sd55;
gen_input_real[819] = -18'sd4;
gen_input_real[115] = 18'sd83;
gen_input_real[371] = 18'sd0;
gen_input_real[627] = -18'sd90;
gen_input_real[883] = -18'sd19;
gen_input_real[179] = 18'sd78;
gen_input_real[435] = 18'sd29;
gen_input_real[691] = -18'sd72;
gen_input_real[947] = -18'sd11;
gen_input_real[243] = 18'sd70;
gen_input_real[499] = -18'sd14;
gen_input_real[755] = -18'sd55;
gen_input_real[1011] = 18'sd29;
gen_input_real[7] = 18'sd27;
gen_input_real[263] = -18'sd33;
gen_input_real[519] = 18'sd8;
gen_input_real[775] = 18'sd29;
gen_input_real[71] = -18'sd41;
gen_input_real[327] = -18'sd11;
gen_input_real[583] = 18'sd52;
gen_input_real[839] = -18'sd14;
gen_input_real[135] = -18'sd34;
gen_input_real[391] = 18'sd15;
gen_input_real[647] = 18'sd16;
gen_input_real[903] = 18'sd3;
gen_input_real[199] = -18'sd28;
gen_input_real[455] = -18'sd15;
gen_input_real[711] = 18'sd52;
gen_input_real[967] = 18'sd24;
gen_input_real[23] = -18'sd55;
gen_input_real[279] = -18'sd31;
gen_input_real[535] = 18'sd36;
gen_input_real[791] = 18'sd27;
gen_input_real[87] = 18'sd0;
gen_input_real[343] = -18'sd24;
gen_input_real[599] = -18'sd41;
gen_input_real[855] = 18'sd21;
gen_input_real[151] = 18'sd46;
gen_input_real[407] = 18'sd14;
gen_input_real[663] = -18'sd12;
gen_input_real[919] = -18'sd85;
gen_input_real[215] = -18'sd12;
gen_input_real[471] = 18'sd124;
gen_input_real[727] = 18'sd5;
gen_input_real[983] = -18'sd89;
gen_input_real[39] = 18'sd19;
gen_input_real[295] = 18'sd26;
gen_input_real[551] = -18'sd34;
gen_input_real[807] = 18'sd10;
gen_input_real[103] = 18'sd29;
gen_input_real[359] = -18'sd24;
gen_input_real[615] = -18'sd15;
gen_input_real[871] = 18'sd32;
gen_input_real[167] = 18'sd5;
gen_input_real[423] = -18'sd36;
gen_input_real[679] = -18'sd2;
gen_input_real[935] = 18'sd30;
gen_input_real[231] = -18'sd2;
gen_input_real[487] = -18'sd20;
gen_input_real[743] = 18'sd12;
gen_input_real[999] = 18'sd29;
gen_input_real[55] = -18'sd19;
gen_input_real[311] = -18'sd58;
gen_input_real[567] = 18'sd18;
gen_input_real[823] = 18'sd90;
gen_input_real[119] = -18'sd3;
gen_input_real[375] = -18'sd109;
gen_input_real[631] = -18'sd21;
gen_input_real[887] = 18'sd102;
gen_input_real[183] = 18'sd35;
gen_input_real[439] = -18'sd72;
gen_input_real[695] = -18'sd24;
gen_input_real[951] = 18'sd42;
gen_input_real[247] = 18'sd0;
gen_input_real[503] = -18'sd29;
gen_input_real[759] = 18'sd23;
gen_input_real[1015] = 18'sd21;
gen_input_real[11] = -18'sd46;
gen_input_real[267] = -18'sd8;
gen_input_real[523] = 18'sd67;
gen_input_real[779] = -18'sd6;
gen_input_real[75] = -18'sd70;
gen_input_real[331] = 18'sd21;
gen_input_real[587] = 18'sd47;
gen_input_real[843] = -18'sd34;
gen_input_real[139] = -18'sd19;
gen_input_real[395] = 18'sd17;
gen_input_real[651] = 18'sd8;
gen_input_real[907] = 18'sd36;
gen_input_real[203] = -18'sd13;
gen_input_real[459] = -18'sd87;
gen_input_real[715] = 18'sd20;
gen_input_real[971] = 18'sd78;
gen_input_real[27] = -18'sd17;
gen_input_real[283] = -18'sd28;
gen_input_real[539] = -18'sd4;
gen_input_real[795] = 18'sd6;
gen_input_real[91] = 18'sd40;
gen_input_real[347] = -18'sd28;
gen_input_real[603] = -18'sd58;
gen_input_real[859] = 18'sd53;
gen_input_real[155] = 18'sd53;
gen_input_real[411] = -18'sd60;
gen_input_real[667] = -18'sd53;
gen_input_real[923] = 18'sd52;
gen_input_real[219] = 18'sd64;
gen_input_real[475] = -18'sd49;
gen_input_real[731] = -18'sd74;
gen_input_real[987] = 18'sd68;
gen_input_real[43] = 18'sd80;
gen_input_real[299] = -18'sd96;
gen_input_real[555] = -18'sd76;
gen_input_real[811] = 18'sd98;
gen_input_real[107] = 18'sd55;
gen_input_real[363] = -18'sd60;
gen_input_real[619] = -18'sd10;
gen_input_real[875] = 18'sd32;
gen_input_real[171] = -18'sd42;
gen_input_real[427] = -18'sd38;
gen_input_real[683] = 18'sd65;
gen_input_real[939] = 18'sd55;
gen_input_real[235] = -18'sd48;
gen_input_real[491] = -18'sd81;
gen_input_real[747] = 18'sd17;
gen_input_real[1003] = 18'sd116;
gen_input_real[59] = 18'sd9;
gen_input_real[315] = -18'sd128;
gen_input_real[571] = -18'sd32;
gen_input_real[827] = 18'sd107;
gen_input_real[123] = 18'sd43;
gen_input_real[379] = -18'sd81;
gen_input_real[635] = -18'sd29;
gen_input_real[891] = 18'sd58;
gen_input_real[187] = 18'sd6;
gen_input_real[443] = -18'sd35;
gen_input_real[699] = -18'sd5;
gen_input_real[955] = 18'sd18;
gen_input_real[251] = 18'sd23;
gen_input_real[507] = -18'sd11;
gen_input_real[763] = -18'sd48;
gen_input_real[1019] = 18'sd9;
gen_input_real[15] = 18'sd75;
gen_input_real[271] = -18'sd11;
gen_input_real[527] = -18'sd88;
gen_input_real[783] = 18'sd17;
gen_input_real[79] = 18'sd93;
gen_input_real[335] = -18'sd12;
gen_input_real[591] = -18'sd104;
gen_input_real[847] = -18'sd4;
gen_input_real[143] = 18'sd105;
gen_input_real[399] = -18'sd2;
gen_input_real[655] = -18'sd77;
gen_input_real[911] = 18'sd39;
gen_input_real[207] = 18'sd32;
gen_input_real[463] = -18'sd72;
gen_input_real[719] = -18'sd14;
gen_input_real[975] = 18'sd76;
gen_input_real[31] = 18'sd44;
gen_input_real[287] = -18'sd70;
gen_input_real[543] = -18'sd89;
gen_input_real[799] = 18'sd77;
gen_input_real[95] = 18'sd104;
gen_input_real[351] = -18'sd90;
gen_input_real[607] = -18'sd91;
gen_input_real[863] = 18'sd101;
gen_input_real[159] = 18'sd93;
gen_input_real[415] = -18'sd107;
gen_input_real[671] = -18'sd115;
gen_input_real[927] = 18'sd103;
gen_input_real[223] = 18'sd120;
gen_input_real[479] = -18'sd87;
gen_input_real[735] = -18'sd92;
gen_input_real[991] = 18'sd67;
gen_input_real[47] = 18'sd56;
gen_input_real[303] = -18'sd36;
gen_input_real[559] = -18'sd30;
gen_input_real[815] = -18'sd6;
gen_input_real[111] = 18'sd20;
gen_input_real[367] = 18'sd31;
gen_input_real[623] = -18'sd34;
gen_input_real[879] = -18'sd16;
gen_input_real[175] = 18'sd65;
gen_input_real[431] = -18'sd11;
gen_input_real[687] = -18'sd75;
gen_input_real[943] = 18'sd22;
gen_input_real[239] = 18'sd52;
gen_input_real[495] = -18'sd9;
gen_input_real[751] = -18'sd40;
gen_input_real[1007] = -18'sd18;
gen_input_real[63] = 18'sd60;
gen_input_real[319] = 18'sd33;
gen_input_real[575] = -18'sd82;
gen_input_real[831] = -18'sd15;
gen_input_real[127] = 18'sd83;
gen_input_real[383] = -18'sd16;
gen_input_real[639] = -18'sd70;
gen_input_real[895] = 18'sd32;
gen_input_real[191] = 18'sd54;
gen_input_real[447] = -18'sd19;
gen_input_real[703] = -18'sd67;
gen_input_real[959] = -18'sd7;
gen_input_real[255] = 18'sd150;
gen_input_real[511] = 18'sd16;
gen_input_real[767] = -18'sd255;
gen_input_real[1023] = 18'sd0;
