0 0
5 -453
22 -902
49 -1350
88 -1805
139 -2273
201 -2733
296 -3439
363 -3686
463 -4183
633 -5135
703 -5183
988 -6663
991 -6162
1174 -6768
1382 -7426
2175 -10936
1752 -8280
2045 -9110
2387 -10052
4414 -17625
2740 -10396
3221 -11639
3801 -13109
8401 -27697
3790 -11964
4528 -13707
5148 -14965
5791 -16185
6501 -17491
7306 -18942
8249 -20628
9405 -22705
10935 -25511
13258 -29909
18183 -39698
78193 -165326
1651 -3383
9613 -19098
14428 -27808
21365 -39971
79227 -143947
11070 -19542
87139 -149514
-4358 7271
7457 -12102
13029 -20576
17611 -27070
22367 -33474
28237 -41158
36967 -52489
55449 -76714
222219 -299628
-19309 25378
14480 -18554
29992 -37474
44078 -53709
61505 -73097
88421 -102505
144614 -163547
506785 -559151
380442 -409538
264420 -277729
-229085 234778
-116220 116220
-76369 74517
-53512 50947
-36979 34352
-22705 20579
-8139 7196
9805 -8458
37678 -31703
100748 -82681
571710 -457566
-263278 205464
-116190 88403
-68806 51030
-28503 20602
144104 -101490
-150328 103136
-89153 59570
-69442 45177
-57635 36497
-48116 29648
-38044 22802
-21826 12720
62810 -35581
-94681 52112
-56033 29950
-37432 19421
22205 -11177
-85122 41545
-56797 26863
-45908 21027
-35177 15593
925 -396
-55213 22870
8296 -3317
-90294 34830
-62854 23363
-54745 19588
-49950 17184
-45591 15061
-33961 10758
-54957 16671
-47808 13864
-45131 12489
-42937 11316
-37944 9504
-46375 11013
-42725 9594
-39553 8373
-43721 8696
-41654 7755
-40726 7066
-39498 6355
-40769 6047
-39882 5416
-39435 4863
-38977 4322
-39109 3851
-38775 3339
-38588 2846
-38415 2360
-38294 1881
-38221 1407
-38153 936
-38120 467
-38112 0
-38120 -467
-38153 -936
-38221 -1407
-38294 -1881
-38415 -2360
-38588 -2846
-38775 -3339
-39109 -3851
-38977 -4322
-39435 -4863
-39882 -5416
-40769 -6047
-39498 -6355
-40726 -7066
-41654 -7755
-43721 -8696
-39553 -8373
-42725 -9594
-46375 -11013
-37944 -9504
-42937 -11316
-45131 -12489
-47808 -13864
-54957 -16671
-33961 -10758
-45591 -15061
-49950 -17184
-54745 -19588
-62854 -23363
-90294 -34830
8296 3317
-55213 -22870
925 396
-35177 -15593
-45908 -21027
-56797 -26863
-85122 -41545
22205 11177
-37432 -19421
-56033 -29950
-94681 -52112
62810 35581
-21826 -12720
-38044 -22802
-48116 -29648
-57635 -36497
-69442 -45177
-89153 -59570
-150328 -103136
144104 101490
-28503 -20602
-68806 -51030
-116190 -88403
-263278 -205464
571710 457566
100748 82681
37678 31703
9805 8458
-8139 -7196
-22705 -20579
-36979 -34352
-53512 -50947
-76369 -74517
-116220 -116220
-229085 -234778
264420 277729
380442 409538
506785 559151
144614 163547
88421 102505
61505 73097
44078 53709
29992 37474
14480 18554
-19309 -25378
222219 299628
55449 76714
36967 52489
28237 41158
22367 33474
17611 27070
13029 20576
7457 12102
-4358 -7271
87139 149514
11070 19542
79227 143947
21365 39971
14428 27808
9613 19098
1651 3383
78193 165326
18183 39698
13258 29909
10935 25511
9405 22705
8249 20628
7306 18942
6501 17491
5791 16185
5148 14965
4528 13707
3790 11964
8401 27697
3801 13109
3221 11639
2740 10396
4414 17625
2387 10052
2045 9110
1752 8280
2175 10936
1382 7426
1174 6768
991 6162
988 6663
703 5183
633 5135
463 4183
363 3686
296 3439
201 2733
139 2273
88 1805
49 1350
22 902
5 453
