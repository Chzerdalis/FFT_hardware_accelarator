w_real[0] = 12'h7FF; w_imag[0] = 12'h000;
w_real[1] = 12'h7FF; w_imag[1] = 12'hFF4;
w_real[2] = 12'h7FF; w_imag[2] = 12'hFE7;
w_real[3] = 12'h7FF; w_imag[3] = 12'hFDB;
w_real[4] = 12'h7FF; w_imag[4] = 12'hFCE;
w_real[5] = 12'h7FF; w_imag[5] = 12'hFC2;
w_real[6] = 12'h7FE; w_imag[6] = 12'hFB5;
w_real[7] = 12'h7FE; w_imag[7] = 12'hFA9;
w_real[8] = 12'h7FD; w_imag[8] = 12'hF9C;
w_real[9] = 12'h7FC; w_imag[9] = 12'hF8F;
w_real[10] = 12'h7FC; w_imag[10] = 12'hF83;
w_real[11] = 12'h7FB; w_imag[11] = 12'hF76;
w_real[12] = 12'h7FA; w_imag[12] = 12'hF6A;
w_real[13] = 12'h7F9; w_imag[13] = 12'hF5D;
w_real[14] = 12'h7F8; w_imag[14] = 12'hF51;
w_real[15] = 12'h7F7; w_imag[15] = 12'hF44;
w_real[16] = 12'h7F6; w_imag[16] = 12'hF38;
w_real[17] = 12'h7F4; w_imag[17] = 12'hF2B;
w_real[18] = 12'h7F3; w_imag[18] = 12'hF1F;
w_real[19] = 12'h7F2; w_imag[19] = 12'hF12;
w_real[20] = 12'h7F0; w_imag[20] = 12'hF06;
w_real[21] = 12'h7EF; w_imag[21] = 12'hEF9;
w_real[22] = 12'h7ED; w_imag[22] = 12'hEED;
w_real[23] = 12'h7EB; w_imag[23] = 12'hEE0;
w_real[24] = 12'h7E9; w_imag[24] = 12'hED4;
w_real[25] = 12'h7E7; w_imag[25] = 12'hEC8;
w_real[26] = 12'h7E5; w_imag[26] = 12'hEBB;
w_real[27] = 12'h7E3; w_imag[27] = 12'hEAF;
w_real[28] = 12'h7E1; w_imag[28] = 12'hEA2;
w_real[29] = 12'h7DF; w_imag[29] = 12'hE96;
w_real[30] = 12'h7DD; w_imag[30] = 12'hE8A;
w_real[31] = 12'h7DB; w_imag[31] = 12'hE7D;
w_real[32] = 12'h7D8; w_imag[32] = 12'hE71;
w_real[33] = 12'h7D6; w_imag[33] = 12'hE65;
w_real[34] = 12'h7D3; w_imag[34] = 12'hE58;
w_real[35] = 12'h7D0; w_imag[35] = 12'hE4C;
w_real[36] = 12'h7CE; w_imag[36] = 12'hE40;
w_real[37] = 12'h7CB; w_imag[37] = 12'hE34;
w_real[38] = 12'h7C8; w_imag[38] = 12'hE27;
w_real[39] = 12'h7C5; w_imag[39] = 12'hE1B;
w_real[40] = 12'h7C2; w_imag[40] = 12'hE0F;
w_real[41] = 12'h7BF; w_imag[41] = 12'hE03;
w_real[42] = 12'h7BC; w_imag[42] = 12'hDF7;
w_real[43] = 12'h7B9; w_imag[43] = 12'hDEA;
w_real[44] = 12'h7B5; w_imag[44] = 12'hDDE;
w_real[45] = 12'h7B2; w_imag[45] = 12'hDD2;
w_real[46] = 12'h7AE; w_imag[46] = 12'hDC6;
w_real[47] = 12'h7AB; w_imag[47] = 12'hDBA;
w_real[48] = 12'h7A7; w_imag[48] = 12'hDAE;
w_real[49] = 12'h7A4; w_imag[49] = 12'hDA2;
w_real[50] = 12'h7A0; w_imag[50] = 12'hD96;
w_real[51] = 12'h79C; w_imag[51] = 12'hD8A;
w_real[52] = 12'h798; w_imag[52] = 12'hD7E;
w_real[53] = 12'h794; w_imag[53] = 12'hD72;
w_real[54] = 12'h790; w_imag[54] = 12'hD66;
w_real[55] = 12'h78C; w_imag[55] = 12'hD5A;
w_real[56] = 12'h788; w_imag[56] = 12'hD4F;
w_real[57] = 12'h784; w_imag[57] = 12'hD43;
w_real[58] = 12'h77F; w_imag[58] = 12'hD37;
w_real[59] = 12'h77B; w_imag[59] = 12'hD2B;
w_real[60] = 12'h776; w_imag[60] = 12'hD1F;
w_real[61] = 12'h772; w_imag[61] = 12'hD14;
w_real[62] = 12'h76D; w_imag[62] = 12'hD08;
w_real[63] = 12'h768; w_imag[63] = 12'hCFC;
w_real[64] = 12'h764; w_imag[64] = 12'hCF1;
w_real[65] = 12'h75F; w_imag[65] = 12'hCE5;
w_real[66] = 12'h75A; w_imag[66] = 12'hCDA;
w_real[67] = 12'h755; w_imag[67] = 12'hCCE;
w_real[68] = 12'h750; w_imag[68] = 12'hCC3;
w_real[69] = 12'h74B; w_imag[69] = 12'hCB7;
w_real[70] = 12'h745; w_imag[70] = 12'hCAC;
w_real[71] = 12'h740; w_imag[71] = 12'hCA0;
w_real[72] = 12'h73B; w_imag[72] = 12'hC95;
w_real[73] = 12'h735; w_imag[73] = 12'hC8A;
w_real[74] = 12'h730; w_imag[74] = 12'hC7E;
w_real[75] = 12'h72A; w_imag[75] = 12'hC73;
w_real[76] = 12'h725; w_imag[76] = 12'hC68;
w_real[77] = 12'h71F; w_imag[77] = 12'hC5C;
w_real[78] = 12'h719; w_imag[78] = 12'hC51;
w_real[79] = 12'h714; w_imag[79] = 12'hC46;
w_real[80] = 12'h70E; w_imag[80] = 12'hC3B;
w_real[81] = 12'h708; w_imag[81] = 12'hC30;
w_real[82] = 12'h702; w_imag[82] = 12'hC25;
w_real[83] = 12'h6FC; w_imag[83] = 12'hC1A;
w_real[84] = 12'h6F5; w_imag[84] = 12'hC0F;
w_real[85] = 12'h6EF; w_imag[85] = 12'hC04;
w_real[86] = 12'h6E9; w_imag[86] = 12'hBF9;
w_real[87] = 12'h6E3; w_imag[87] = 12'hBEE;
w_real[88] = 12'h6DC; w_imag[88] = 12'hBE4;
w_real[89] = 12'h6D6; w_imag[89] = 12'hBD9;
w_real[90] = 12'h6CF; w_imag[90] = 12'hBCE;
w_real[91] = 12'h6C8; w_imag[91] = 12'hBC3;
w_real[92] = 12'h6C2; w_imag[92] = 12'hBB9;
w_real[93] = 12'h6BB; w_imag[93] = 12'hBAE;
w_real[94] = 12'h6B4; w_imag[94] = 12'hBA4;
w_real[95] = 12'h6AD; w_imag[95] = 12'hB99;
w_real[96] = 12'h6A6; w_imag[96] = 12'hB8F;
w_real[97] = 12'h69F; w_imag[97] = 12'hB84;
w_real[98] = 12'h698; w_imag[98] = 12'hB7A;
w_real[99] = 12'h691; w_imag[99] = 12'hB70;
w_real[100] = 12'h68A; w_imag[100] = 12'hB65;
w_real[101] = 12'h683; w_imag[101] = 12'hB5B;
w_real[102] = 12'h67B; w_imag[102] = 12'hB51;
w_real[103] = 12'h674; w_imag[103] = 12'hB47;
w_real[104] = 12'h66C; w_imag[104] = 12'hB3D;
w_real[105] = 12'h665; w_imag[105] = 12'hB32;
w_real[106] = 12'h65D; w_imag[106] = 12'hB28;
w_real[107] = 12'h656; w_imag[107] = 12'hB1E;
w_real[108] = 12'h64E; w_imag[108] = 12'hB15;
w_real[109] = 12'h646; w_imag[109] = 12'hB0B;
w_real[110] = 12'h63E; w_imag[110] = 12'hB01;
w_real[111] = 12'h637; w_imag[111] = 12'hAF7;
w_real[112] = 12'h62F; w_imag[112] = 12'hAED;
w_real[113] = 12'h627; w_imag[113] = 12'hAE4;
w_real[114] = 12'h61F; w_imag[114] = 12'hADA;
w_real[115] = 12'h616; w_imag[115] = 12'hAD0;
w_real[116] = 12'h60E; w_imag[116] = 12'hAC7;
w_real[117] = 12'h606; w_imag[117] = 12'hABD;
w_real[118] = 12'h5FE; w_imag[118] = 12'hAB4;
w_real[119] = 12'h5F5; w_imag[119] = 12'hAAA;
w_real[120] = 12'h5ED; w_imag[120] = 12'hAA1;
w_real[121] = 12'h5E5; w_imag[121] = 12'hA98;
w_real[122] = 12'h5DC; w_imag[122] = 12'hA8F;
w_real[123] = 12'h5D3; w_imag[123] = 12'hA85;
w_real[124] = 12'h5CB; w_imag[124] = 12'hA7C;
w_real[125] = 12'h5C2; w_imag[125] = 12'hA73;
w_real[126] = 12'h5B9; w_imag[126] = 12'hA6A;
w_real[127] = 12'h5B1; w_imag[127] = 12'hA61;
w_real[128] = 12'h5A8; w_imag[128] = 12'hA58;
w_real[129] = 12'h59F; w_imag[129] = 12'hA4F;
w_real[130] = 12'h596; w_imag[130] = 12'hA47;
w_real[131] = 12'h58D; w_imag[131] = 12'hA3E;
w_real[132] = 12'h584; w_imag[132] = 12'hA35;
w_real[133] = 12'h57B; w_imag[133] = 12'hA2D;
w_real[134] = 12'h571; w_imag[134] = 12'hA24;
w_real[135] = 12'h568; w_imag[135] = 12'hA1B;
w_real[136] = 12'h55F; w_imag[136] = 12'hA13;
w_real[137] = 12'h556; w_imag[137] = 12'hA0B;
w_real[138] = 12'h54C; w_imag[138] = 12'hA02;
w_real[139] = 12'h543; w_imag[139] = 12'h9FA;
w_real[140] = 12'h539; w_imag[140] = 12'h9F2;
w_real[141] = 12'h530; w_imag[141] = 12'h9EA;
w_real[142] = 12'h526; w_imag[142] = 12'h9E1;
w_real[143] = 12'h51C; w_imag[143] = 12'h9D9;
w_real[144] = 12'h513; w_imag[144] = 12'h9D1;
w_real[145] = 12'h509; w_imag[145] = 12'h9C9;
w_real[146] = 12'h4FF; w_imag[146] = 12'h9C2;
w_real[147] = 12'h4F5; w_imag[147] = 12'h9BA;
w_real[148] = 12'h4EB; w_imag[148] = 12'h9B2;
w_real[149] = 12'h4E2; w_imag[149] = 12'h9AA;
w_real[150] = 12'h4D8; w_imag[150] = 12'h9A3;
w_real[151] = 12'h4CE; w_imag[151] = 12'h99B;
w_real[152] = 12'h4C3; w_imag[152] = 12'h994;
w_real[153] = 12'h4B9; w_imag[153] = 12'h98C;
w_real[154] = 12'h4AF; w_imag[154] = 12'h985;
w_real[155] = 12'h4A5; w_imag[155] = 12'h97D;
w_real[156] = 12'h49B; w_imag[156] = 12'h976;
w_real[157] = 12'h490; w_imag[157] = 12'h96F;
w_real[158] = 12'h486; w_imag[158] = 12'h968;
w_real[159] = 12'h47C; w_imag[159] = 12'h961;
w_real[160] = 12'h471; w_imag[160] = 12'h95A;
w_real[161] = 12'h467; w_imag[161] = 12'h953;
w_real[162] = 12'h45C; w_imag[162] = 12'h94C;
w_real[163] = 12'h452; w_imag[163] = 12'h945;
w_real[164] = 12'h447; w_imag[164] = 12'h93E;
w_real[165] = 12'h43D; w_imag[165] = 12'h938;
w_real[166] = 12'h432; w_imag[166] = 12'h931;
w_real[167] = 12'h427; w_imag[167] = 12'h92A;
w_real[168] = 12'h41C; w_imag[168] = 12'h924;
w_real[169] = 12'h412; w_imag[169] = 12'h91D;
w_real[170] = 12'h407; w_imag[170] = 12'h917;
w_real[171] = 12'h3FC; w_imag[171] = 12'h911;
w_real[172] = 12'h3F1; w_imag[172] = 12'h90B;
w_real[173] = 12'h3E6; w_imag[173] = 12'h904;
w_real[174] = 12'h3DB; w_imag[174] = 12'h8FE;
w_real[175] = 12'h3D0; w_imag[175] = 12'h8F8;
w_real[176] = 12'h3C5; w_imag[176] = 12'h8F2;
w_real[177] = 12'h3BA; w_imag[177] = 12'h8EC;
w_real[178] = 12'h3AF; w_imag[178] = 12'h8E7;
w_real[179] = 12'h3A4; w_imag[179] = 12'h8E1;
w_real[180] = 12'h398; w_imag[180] = 12'h8DB;
w_real[181] = 12'h38D; w_imag[181] = 12'h8D6;
w_real[182] = 12'h382; w_imag[182] = 12'h8D0;
w_real[183] = 12'h376; w_imag[183] = 12'h8CB;
w_real[184] = 12'h36B; w_imag[184] = 12'h8C5;
w_real[185] = 12'h360; w_imag[185] = 12'h8C0;
w_real[186] = 12'h354; w_imag[186] = 12'h8BB;
w_real[187] = 12'h349; w_imag[187] = 12'h8B5;
w_real[188] = 12'h33D; w_imag[188] = 12'h8B0;
w_real[189] = 12'h332; w_imag[189] = 12'h8AB;
w_real[190] = 12'h326; w_imag[190] = 12'h8A6;
w_real[191] = 12'h31B; w_imag[191] = 12'h8A1;
w_real[192] = 12'h30F; w_imag[192] = 12'h89C;
w_real[193] = 12'h304; w_imag[193] = 12'h898;
w_real[194] = 12'h2F8; w_imag[194] = 12'h893;
w_real[195] = 12'h2EC; w_imag[195] = 12'h88E;
w_real[196] = 12'h2E1; w_imag[196] = 12'h88A;
w_real[197] = 12'h2D5; w_imag[197] = 12'h885;
w_real[198] = 12'h2C9; w_imag[198] = 12'h881;
w_real[199] = 12'h2BD; w_imag[199] = 12'h87C;
w_real[200] = 12'h2B1; w_imag[200] = 12'h878;
w_real[201] = 12'h2A6; w_imag[201] = 12'h874;
w_real[202] = 12'h29A; w_imag[202] = 12'h870;
w_real[203] = 12'h28E; w_imag[203] = 12'h86C;
w_real[204] = 12'h282; w_imag[204] = 12'h868;
w_real[205] = 12'h276; w_imag[205] = 12'h864;
w_real[206] = 12'h26A; w_imag[206] = 12'h860;
w_real[207] = 12'h25E; w_imag[207] = 12'h85C;
w_real[208] = 12'h252; w_imag[208] = 12'h859;
w_real[209] = 12'h246; w_imag[209] = 12'h855;
w_real[210] = 12'h23A; w_imag[210] = 12'h852;
w_real[211] = 12'h22E; w_imag[211] = 12'h84E;
w_real[212] = 12'h222; w_imag[212] = 12'h84B;
w_real[213] = 12'h216; w_imag[213] = 12'h847;
w_real[214] = 12'h209; w_imag[214] = 12'h844;
w_real[215] = 12'h1FD; w_imag[215] = 12'h841;
w_real[216] = 12'h1F1; w_imag[216] = 12'h83E;
w_real[217] = 12'h1E5; w_imag[217] = 12'h83B;
w_real[218] = 12'h1D9; w_imag[218] = 12'h838;
w_real[219] = 12'h1CC; w_imag[219] = 12'h835;
w_real[220] = 12'h1C0; w_imag[220] = 12'h832;
w_real[221] = 12'h1B4; w_imag[221] = 12'h830;
w_real[222] = 12'h1A8; w_imag[222] = 12'h82D;
w_real[223] = 12'h19B; w_imag[223] = 12'h82A;
w_real[224] = 12'h18F; w_imag[224] = 12'h828;
w_real[225] = 12'h183; w_imag[225] = 12'h825;
w_real[226] = 12'h176; w_imag[226] = 12'h823;
w_real[227] = 12'h16A; w_imag[227] = 12'h821;
w_real[228] = 12'h15E; w_imag[228] = 12'h81F;
w_real[229] = 12'h151; w_imag[229] = 12'h81D;
w_real[230] = 12'h145; w_imag[230] = 12'h81B;
w_real[231] = 12'h138; w_imag[231] = 12'h819;
w_real[232] = 12'h12C; w_imag[232] = 12'h817;
w_real[233] = 12'h120; w_imag[233] = 12'h815;
w_real[234] = 12'h113; w_imag[234] = 12'h813;
w_real[235] = 12'h107; w_imag[235] = 12'h811;
w_real[236] = 12'h0FA; w_imag[236] = 12'h810;
w_real[237] = 12'h0EE; w_imag[237] = 12'h80E;
w_real[238] = 12'h0E1; w_imag[238] = 12'h80D;
w_real[239] = 12'h0D5; w_imag[239] = 12'h80C;
w_real[240] = 12'h0C8; w_imag[240] = 12'h80A;
w_real[241] = 12'h0BC; w_imag[241] = 12'h809;
w_real[242] = 12'h0AF; w_imag[242] = 12'h808;
w_real[243] = 12'h0A3; w_imag[243] = 12'h807;
w_real[244] = 12'h096; w_imag[244] = 12'h806;
w_real[245] = 12'h08A; w_imag[245] = 12'h805;
w_real[246] = 12'h07D; w_imag[246] = 12'h804;
w_real[247] = 12'h071; w_imag[247] = 12'h804;
w_real[248] = 12'h064; w_imag[248] = 12'h803;
w_real[249] = 12'h057; w_imag[249] = 12'h802;
w_real[250] = 12'h04B; w_imag[250] = 12'h802;
w_real[251] = 12'h03E; w_imag[251] = 12'h801;
w_real[252] = 12'h032; w_imag[252] = 12'h801;
w_real[253] = 12'h025; w_imag[253] = 12'h801;
w_real[254] = 12'h019; w_imag[254] = 12'h801;
w_real[255] = 12'h00C; w_imag[255] = 12'h801;
w_real[256] = 12'h000; w_imag[256] = 12'h800;
w_real[257] = 12'hFF4; w_imag[257] = 12'h801;
w_real[258] = 12'hFE7; w_imag[258] = 12'h801;
w_real[259] = 12'hFDB; w_imag[259] = 12'h801;
w_real[260] = 12'hFCE; w_imag[260] = 12'h801;
w_real[261] = 12'hFC2; w_imag[261] = 12'h801;
w_real[262] = 12'hFB5; w_imag[262] = 12'h802;
w_real[263] = 12'hFA9; w_imag[263] = 12'h802;
w_real[264] = 12'hF9C; w_imag[264] = 12'h803;
w_real[265] = 12'hF8F; w_imag[265] = 12'h804;
w_real[266] = 12'hF83; w_imag[266] = 12'h804;
w_real[267] = 12'hF76; w_imag[267] = 12'h805;
w_real[268] = 12'hF6A; w_imag[268] = 12'h806;
w_real[269] = 12'hF5D; w_imag[269] = 12'h807;
w_real[270] = 12'hF51; w_imag[270] = 12'h808;
w_real[271] = 12'hF44; w_imag[271] = 12'h809;
w_real[272] = 12'hF38; w_imag[272] = 12'h80A;
w_real[273] = 12'hF2B; w_imag[273] = 12'h80C;
w_real[274] = 12'hF1F; w_imag[274] = 12'h80D;
w_real[275] = 12'hF12; w_imag[275] = 12'h80E;
w_real[276] = 12'hF06; w_imag[276] = 12'h810;
w_real[277] = 12'hEF9; w_imag[277] = 12'h811;
w_real[278] = 12'hEED; w_imag[278] = 12'h813;
w_real[279] = 12'hEE0; w_imag[279] = 12'h815;
w_real[280] = 12'hED4; w_imag[280] = 12'h817;
w_real[281] = 12'hEC8; w_imag[281] = 12'h819;
w_real[282] = 12'hEBB; w_imag[282] = 12'h81B;
w_real[283] = 12'hEAF; w_imag[283] = 12'h81D;
w_real[284] = 12'hEA2; w_imag[284] = 12'h81F;
w_real[285] = 12'hE96; w_imag[285] = 12'h821;
w_real[286] = 12'hE8A; w_imag[286] = 12'h823;
w_real[287] = 12'hE7D; w_imag[287] = 12'h825;
w_real[288] = 12'hE71; w_imag[288] = 12'h828;
w_real[289] = 12'hE65; w_imag[289] = 12'h82A;
w_real[290] = 12'hE58; w_imag[290] = 12'h82D;
w_real[291] = 12'hE4C; w_imag[291] = 12'h830;
w_real[292] = 12'hE40; w_imag[292] = 12'h832;
w_real[293] = 12'hE34; w_imag[293] = 12'h835;
w_real[294] = 12'hE27; w_imag[294] = 12'h838;
w_real[295] = 12'hE1B; w_imag[295] = 12'h83B;
w_real[296] = 12'hE0F; w_imag[296] = 12'h83E;
w_real[297] = 12'hE03; w_imag[297] = 12'h841;
w_real[298] = 12'hDF7; w_imag[298] = 12'h844;
w_real[299] = 12'hDEA; w_imag[299] = 12'h847;
w_real[300] = 12'hDDE; w_imag[300] = 12'h84B;
w_real[301] = 12'hDD2; w_imag[301] = 12'h84E;
w_real[302] = 12'hDC6; w_imag[302] = 12'h852;
w_real[303] = 12'hDBA; w_imag[303] = 12'h855;
w_real[304] = 12'hDAE; w_imag[304] = 12'h859;
w_real[305] = 12'hDA2; w_imag[305] = 12'h85C;
w_real[306] = 12'hD96; w_imag[306] = 12'h860;
w_real[307] = 12'hD8A; w_imag[307] = 12'h864;
w_real[308] = 12'hD7E; w_imag[308] = 12'h868;
w_real[309] = 12'hD72; w_imag[309] = 12'h86C;
w_real[310] = 12'hD66; w_imag[310] = 12'h870;
w_real[311] = 12'hD5A; w_imag[311] = 12'h874;
w_real[312] = 12'hD4F; w_imag[312] = 12'h878;
w_real[313] = 12'hD43; w_imag[313] = 12'h87C;
w_real[314] = 12'hD37; w_imag[314] = 12'h881;
w_real[315] = 12'hD2B; w_imag[315] = 12'h885;
w_real[316] = 12'hD1F; w_imag[316] = 12'h88A;
w_real[317] = 12'hD14; w_imag[317] = 12'h88E;
w_real[318] = 12'hD08; w_imag[318] = 12'h893;
w_real[319] = 12'hCFC; w_imag[319] = 12'h898;
w_real[320] = 12'hCF1; w_imag[320] = 12'h89C;
w_real[321] = 12'hCE5; w_imag[321] = 12'h8A1;
w_real[322] = 12'hCDA; w_imag[322] = 12'h8A6;
w_real[323] = 12'hCCE; w_imag[323] = 12'h8AB;
w_real[324] = 12'hCC3; w_imag[324] = 12'h8B0;
w_real[325] = 12'hCB7; w_imag[325] = 12'h8B5;
w_real[326] = 12'hCAC; w_imag[326] = 12'h8BB;
w_real[327] = 12'hCA0; w_imag[327] = 12'h8C0;
w_real[328] = 12'hC95; w_imag[328] = 12'h8C5;
w_real[329] = 12'hC8A; w_imag[329] = 12'h8CB;
w_real[330] = 12'hC7E; w_imag[330] = 12'h8D0;
w_real[331] = 12'hC73; w_imag[331] = 12'h8D6;
w_real[332] = 12'hC68; w_imag[332] = 12'h8DB;
w_real[333] = 12'hC5C; w_imag[333] = 12'h8E1;
w_real[334] = 12'hC51; w_imag[334] = 12'h8E7;
w_real[335] = 12'hC46; w_imag[335] = 12'h8EC;
w_real[336] = 12'hC3B; w_imag[336] = 12'h8F2;
w_real[337] = 12'hC30; w_imag[337] = 12'h8F8;
w_real[338] = 12'hC25; w_imag[338] = 12'h8FE;
w_real[339] = 12'hC1A; w_imag[339] = 12'h904;
w_real[340] = 12'hC0F; w_imag[340] = 12'h90B;
w_real[341] = 12'hC04; w_imag[341] = 12'h911;
w_real[342] = 12'hBF9; w_imag[342] = 12'h917;
w_real[343] = 12'hBEE; w_imag[343] = 12'h91D;
w_real[344] = 12'hBE4; w_imag[344] = 12'h924;
w_real[345] = 12'hBD9; w_imag[345] = 12'h92A;
w_real[346] = 12'hBCE; w_imag[346] = 12'h931;
w_real[347] = 12'hBC3; w_imag[347] = 12'h938;
w_real[348] = 12'hBB9; w_imag[348] = 12'h93E;
w_real[349] = 12'hBAE; w_imag[349] = 12'h945;
w_real[350] = 12'hBA4; w_imag[350] = 12'h94C;
w_real[351] = 12'hB99; w_imag[351] = 12'h953;
w_real[352] = 12'hB8F; w_imag[352] = 12'h95A;
w_real[353] = 12'hB84; w_imag[353] = 12'h961;
w_real[354] = 12'hB7A; w_imag[354] = 12'h968;
w_real[355] = 12'hB70; w_imag[355] = 12'h96F;
w_real[356] = 12'hB65; w_imag[356] = 12'h976;
w_real[357] = 12'hB5B; w_imag[357] = 12'h97D;
w_real[358] = 12'hB51; w_imag[358] = 12'h985;
w_real[359] = 12'hB47; w_imag[359] = 12'h98C;
w_real[360] = 12'hB3D; w_imag[360] = 12'h994;
w_real[361] = 12'hB32; w_imag[361] = 12'h99B;
w_real[362] = 12'hB28; w_imag[362] = 12'h9A3;
w_real[363] = 12'hB1E; w_imag[363] = 12'h9AA;
w_real[364] = 12'hB15; w_imag[364] = 12'h9B2;
w_real[365] = 12'hB0B; w_imag[365] = 12'h9BA;
w_real[366] = 12'hB01; w_imag[366] = 12'h9C2;
w_real[367] = 12'hAF7; w_imag[367] = 12'h9C9;
w_real[368] = 12'hAED; w_imag[368] = 12'h9D1;
w_real[369] = 12'hAE4; w_imag[369] = 12'h9D9;
w_real[370] = 12'hADA; w_imag[370] = 12'h9E1;
w_real[371] = 12'hAD0; w_imag[371] = 12'h9EA;
w_real[372] = 12'hAC7; w_imag[372] = 12'h9F2;
w_real[373] = 12'hABD; w_imag[373] = 12'h9FA;
w_real[374] = 12'hAB4; w_imag[374] = 12'hA02;
w_real[375] = 12'hAAA; w_imag[375] = 12'hA0B;
w_real[376] = 12'hAA1; w_imag[376] = 12'hA13;
w_real[377] = 12'hA98; w_imag[377] = 12'hA1B;
w_real[378] = 12'hA8F; w_imag[378] = 12'hA24;
w_real[379] = 12'hA85; w_imag[379] = 12'hA2D;
w_real[380] = 12'hA7C; w_imag[380] = 12'hA35;
w_real[381] = 12'hA73; w_imag[381] = 12'hA3E;
w_real[382] = 12'hA6A; w_imag[382] = 12'hA47;
w_real[383] = 12'hA61; w_imag[383] = 12'hA4F;
w_real[384] = 12'hA58; w_imag[384] = 12'hA58;
w_real[385] = 12'hA4F; w_imag[385] = 12'hA61;
w_real[386] = 12'hA47; w_imag[386] = 12'hA6A;
w_real[387] = 12'hA3E; w_imag[387] = 12'hA73;
w_real[388] = 12'hA35; w_imag[388] = 12'hA7C;
w_real[389] = 12'hA2D; w_imag[389] = 12'hA85;
w_real[390] = 12'hA24; w_imag[390] = 12'hA8F;
w_real[391] = 12'hA1B; w_imag[391] = 12'hA98;
w_real[392] = 12'hA13; w_imag[392] = 12'hAA1;
w_real[393] = 12'hA0B; w_imag[393] = 12'hAAA;
w_real[394] = 12'hA02; w_imag[394] = 12'hAB4;
w_real[395] = 12'h9FA; w_imag[395] = 12'hABD;
w_real[396] = 12'h9F2; w_imag[396] = 12'hAC7;
w_real[397] = 12'h9EA; w_imag[397] = 12'hAD0;
w_real[398] = 12'h9E1; w_imag[398] = 12'hADA;
w_real[399] = 12'h9D9; w_imag[399] = 12'hAE4;
w_real[400] = 12'h9D1; w_imag[400] = 12'hAED;
w_real[401] = 12'h9C9; w_imag[401] = 12'hAF7;
w_real[402] = 12'h9C2; w_imag[402] = 12'hB01;
w_real[403] = 12'h9BA; w_imag[403] = 12'hB0B;
w_real[404] = 12'h9B2; w_imag[404] = 12'hB15;
w_real[405] = 12'h9AA; w_imag[405] = 12'hB1E;
w_real[406] = 12'h9A3; w_imag[406] = 12'hB28;
w_real[407] = 12'h99B; w_imag[407] = 12'hB32;
w_real[408] = 12'h994; w_imag[408] = 12'hB3D;
w_real[409] = 12'h98C; w_imag[409] = 12'hB47;
w_real[410] = 12'h985; w_imag[410] = 12'hB51;
w_real[411] = 12'h97D; w_imag[411] = 12'hB5B;
w_real[412] = 12'h976; w_imag[412] = 12'hB65;
w_real[413] = 12'h96F; w_imag[413] = 12'hB70;
w_real[414] = 12'h968; w_imag[414] = 12'hB7A;
w_real[415] = 12'h961; w_imag[415] = 12'hB84;
w_real[416] = 12'h95A; w_imag[416] = 12'hB8F;
w_real[417] = 12'h953; w_imag[417] = 12'hB99;
w_real[418] = 12'h94C; w_imag[418] = 12'hBA4;
w_real[419] = 12'h945; w_imag[419] = 12'hBAE;
w_real[420] = 12'h93E; w_imag[420] = 12'hBB9;
w_real[421] = 12'h938; w_imag[421] = 12'hBC3;
w_real[422] = 12'h931; w_imag[422] = 12'hBCE;
w_real[423] = 12'h92A; w_imag[423] = 12'hBD9;
w_real[424] = 12'h924; w_imag[424] = 12'hBE4;
w_real[425] = 12'h91D; w_imag[425] = 12'hBEE;
w_real[426] = 12'h917; w_imag[426] = 12'hBF9;
w_real[427] = 12'h911; w_imag[427] = 12'hC04;
w_real[428] = 12'h90B; w_imag[428] = 12'hC0F;
w_real[429] = 12'h904; w_imag[429] = 12'hC1A;
w_real[430] = 12'h8FE; w_imag[430] = 12'hC25;
w_real[431] = 12'h8F8; w_imag[431] = 12'hC30;
w_real[432] = 12'h8F2; w_imag[432] = 12'hC3B;
w_real[433] = 12'h8EC; w_imag[433] = 12'hC46;
w_real[434] = 12'h8E7; w_imag[434] = 12'hC51;
w_real[435] = 12'h8E1; w_imag[435] = 12'hC5C;
w_real[436] = 12'h8DB; w_imag[436] = 12'hC68;
w_real[437] = 12'h8D6; w_imag[437] = 12'hC73;
w_real[438] = 12'h8D0; w_imag[438] = 12'hC7E;
w_real[439] = 12'h8CB; w_imag[439] = 12'hC8A;
w_real[440] = 12'h8C5; w_imag[440] = 12'hC95;
w_real[441] = 12'h8C0; w_imag[441] = 12'hCA0;
w_real[442] = 12'h8BB; w_imag[442] = 12'hCAC;
w_real[443] = 12'h8B5; w_imag[443] = 12'hCB7;
w_real[444] = 12'h8B0; w_imag[444] = 12'hCC3;
w_real[445] = 12'h8AB; w_imag[445] = 12'hCCE;
w_real[446] = 12'h8A6; w_imag[446] = 12'hCDA;
w_real[447] = 12'h8A1; w_imag[447] = 12'hCE5;
w_real[448] = 12'h89C; w_imag[448] = 12'hCF1;
w_real[449] = 12'h898; w_imag[449] = 12'hCFC;
w_real[450] = 12'h893; w_imag[450] = 12'hD08;
w_real[451] = 12'h88E; w_imag[451] = 12'hD14;
w_real[452] = 12'h88A; w_imag[452] = 12'hD1F;
w_real[453] = 12'h885; w_imag[453] = 12'hD2B;
w_real[454] = 12'h881; w_imag[454] = 12'hD37;
w_real[455] = 12'h87C; w_imag[455] = 12'hD43;
w_real[456] = 12'h878; w_imag[456] = 12'hD4F;
w_real[457] = 12'h874; w_imag[457] = 12'hD5A;
w_real[458] = 12'h870; w_imag[458] = 12'hD66;
w_real[459] = 12'h86C; w_imag[459] = 12'hD72;
w_real[460] = 12'h868; w_imag[460] = 12'hD7E;
w_real[461] = 12'h864; w_imag[461] = 12'hD8A;
w_real[462] = 12'h860; w_imag[462] = 12'hD96;
w_real[463] = 12'h85C; w_imag[463] = 12'hDA2;
w_real[464] = 12'h859; w_imag[464] = 12'hDAE;
w_real[465] = 12'h855; w_imag[465] = 12'hDBA;
w_real[466] = 12'h852; w_imag[466] = 12'hDC6;
w_real[467] = 12'h84E; w_imag[467] = 12'hDD2;
w_real[468] = 12'h84B; w_imag[468] = 12'hDDE;
w_real[469] = 12'h847; w_imag[469] = 12'hDEA;
w_real[470] = 12'h844; w_imag[470] = 12'hDF7;
w_real[471] = 12'h841; w_imag[471] = 12'hE03;
w_real[472] = 12'h83E; w_imag[472] = 12'hE0F;
w_real[473] = 12'h83B; w_imag[473] = 12'hE1B;
w_real[474] = 12'h838; w_imag[474] = 12'hE27;
w_real[475] = 12'h835; w_imag[475] = 12'hE34;
w_real[476] = 12'h832; w_imag[476] = 12'hE40;
w_real[477] = 12'h830; w_imag[477] = 12'hE4C;
w_real[478] = 12'h82D; w_imag[478] = 12'hE58;
w_real[479] = 12'h82A; w_imag[479] = 12'hE65;
w_real[480] = 12'h828; w_imag[480] = 12'hE71;
w_real[481] = 12'h825; w_imag[481] = 12'hE7D;
w_real[482] = 12'h823; w_imag[482] = 12'hE8A;
w_real[483] = 12'h821; w_imag[483] = 12'hE96;
w_real[484] = 12'h81F; w_imag[484] = 12'hEA2;
w_real[485] = 12'h81D; w_imag[485] = 12'hEAF;
w_real[486] = 12'h81B; w_imag[486] = 12'hEBB;
w_real[487] = 12'h819; w_imag[487] = 12'hEC8;
w_real[488] = 12'h817; w_imag[488] = 12'hED4;
w_real[489] = 12'h815; w_imag[489] = 12'hEE0;
w_real[490] = 12'h813; w_imag[490] = 12'hEED;
w_real[491] = 12'h811; w_imag[491] = 12'hEF9;
w_real[492] = 12'h810; w_imag[492] = 12'hF06;
w_real[493] = 12'h80E; w_imag[493] = 12'hF12;
w_real[494] = 12'h80D; w_imag[494] = 12'hF1F;
w_real[495] = 12'h80C; w_imag[495] = 12'hF2B;
w_real[496] = 12'h80A; w_imag[496] = 12'hF38;
w_real[497] = 12'h809; w_imag[497] = 12'hF44;
w_real[498] = 12'h808; w_imag[498] = 12'hF51;
w_real[499] = 12'h807; w_imag[499] = 12'hF5D;
w_real[500] = 12'h806; w_imag[500] = 12'hF6A;
w_real[501] = 12'h805; w_imag[501] = 12'hF76;
w_real[502] = 12'h804; w_imag[502] = 12'hF83;
w_real[503] = 12'h804; w_imag[503] = 12'hF8F;
w_real[504] = 12'h803; w_imag[504] = 12'hF9C;
w_real[505] = 12'h802; w_imag[505] = 12'hFA9;
w_real[506] = 12'h802; w_imag[506] = 12'hFB5;
w_real[507] = 12'h801; w_imag[507] = 12'hFC2;
w_real[508] = 12'h801; w_imag[508] = 12'hFCE;
w_real[509] = 12'h801; w_imag[509] = 12'hFDB;
w_real[510] = 12'h801; w_imag[510] = 12'hFE7;
w_real[511] = 12'h801; w_imag[511] = 12'hFF4;
w_real[512] = 12'h800; w_imag[512] = 12'h000;
w_real[513] = 12'h801; w_imag[513] = 12'h00C;
w_real[514] = 12'h801; w_imag[514] = 12'h019;
w_real[515] = 12'h801; w_imag[515] = 12'h025;
w_real[516] = 12'h801; w_imag[516] = 12'h032;
w_real[517] = 12'h801; w_imag[517] = 12'h03E;
w_real[518] = 12'h802; w_imag[518] = 12'h04B;
w_real[519] = 12'h802; w_imag[519] = 12'h057;
w_real[520] = 12'h803; w_imag[520] = 12'h064;
w_real[521] = 12'h804; w_imag[521] = 12'h071;
w_real[522] = 12'h804; w_imag[522] = 12'h07D;
w_real[523] = 12'h805; w_imag[523] = 12'h08A;
w_real[524] = 12'h806; w_imag[524] = 12'h096;
w_real[525] = 12'h807; w_imag[525] = 12'h0A3;
w_real[526] = 12'h808; w_imag[526] = 12'h0AF;
w_real[527] = 12'h809; w_imag[527] = 12'h0BC;
w_real[528] = 12'h80A; w_imag[528] = 12'h0C8;
w_real[529] = 12'h80C; w_imag[529] = 12'h0D5;
w_real[530] = 12'h80D; w_imag[530] = 12'h0E1;
w_real[531] = 12'h80E; w_imag[531] = 12'h0EE;
w_real[532] = 12'h810; w_imag[532] = 12'h0FA;
w_real[533] = 12'h811; w_imag[533] = 12'h107;
w_real[534] = 12'h813; w_imag[534] = 12'h113;
w_real[535] = 12'h815; w_imag[535] = 12'h120;
w_real[536] = 12'h817; w_imag[536] = 12'h12C;
w_real[537] = 12'h819; w_imag[537] = 12'h138;
w_real[538] = 12'h81B; w_imag[538] = 12'h145;
w_real[539] = 12'h81D; w_imag[539] = 12'h151;
w_real[540] = 12'h81F; w_imag[540] = 12'h15E;
w_real[541] = 12'h821; w_imag[541] = 12'h16A;
w_real[542] = 12'h823; w_imag[542] = 12'h176;
w_real[543] = 12'h825; w_imag[543] = 12'h183;
w_real[544] = 12'h828; w_imag[544] = 12'h18F;
w_real[545] = 12'h82A; w_imag[545] = 12'h19B;
w_real[546] = 12'h82D; w_imag[546] = 12'h1A8;
w_real[547] = 12'h830; w_imag[547] = 12'h1B4;
w_real[548] = 12'h832; w_imag[548] = 12'h1C0;
w_real[549] = 12'h835; w_imag[549] = 12'h1CC;
w_real[550] = 12'h838; w_imag[550] = 12'h1D9;
w_real[551] = 12'h83B; w_imag[551] = 12'h1E5;
w_real[552] = 12'h83E; w_imag[552] = 12'h1F1;
w_real[553] = 12'h841; w_imag[553] = 12'h1FD;
w_real[554] = 12'h844; w_imag[554] = 12'h209;
w_real[555] = 12'h847; w_imag[555] = 12'h216;
w_real[556] = 12'h84B; w_imag[556] = 12'h222;
w_real[557] = 12'h84E; w_imag[557] = 12'h22E;
w_real[558] = 12'h852; w_imag[558] = 12'h23A;
w_real[559] = 12'h855; w_imag[559] = 12'h246;
w_real[560] = 12'h859; w_imag[560] = 12'h252;
w_real[561] = 12'h85C; w_imag[561] = 12'h25E;
w_real[562] = 12'h860; w_imag[562] = 12'h26A;
w_real[563] = 12'h864; w_imag[563] = 12'h276;
w_real[564] = 12'h868; w_imag[564] = 12'h282;
w_real[565] = 12'h86C; w_imag[565] = 12'h28E;
w_real[566] = 12'h870; w_imag[566] = 12'h29A;
w_real[567] = 12'h874; w_imag[567] = 12'h2A6;
w_real[568] = 12'h878; w_imag[568] = 12'h2B1;
w_real[569] = 12'h87C; w_imag[569] = 12'h2BD;
w_real[570] = 12'h881; w_imag[570] = 12'h2C9;
w_real[571] = 12'h885; w_imag[571] = 12'h2D5;
w_real[572] = 12'h88A; w_imag[572] = 12'h2E1;
w_real[573] = 12'h88E; w_imag[573] = 12'h2EC;
w_real[574] = 12'h893; w_imag[574] = 12'h2F8;
w_real[575] = 12'h898; w_imag[575] = 12'h304;
w_real[576] = 12'h89C; w_imag[576] = 12'h30F;
w_real[577] = 12'h8A1; w_imag[577] = 12'h31B;
w_real[578] = 12'h8A6; w_imag[578] = 12'h326;
w_real[579] = 12'h8AB; w_imag[579] = 12'h332;
w_real[580] = 12'h8B0; w_imag[580] = 12'h33D;
w_real[581] = 12'h8B5; w_imag[581] = 12'h349;
w_real[582] = 12'h8BB; w_imag[582] = 12'h354;
w_real[583] = 12'h8C0; w_imag[583] = 12'h360;
w_real[584] = 12'h8C5; w_imag[584] = 12'h36B;
w_real[585] = 12'h8CB; w_imag[585] = 12'h376;
w_real[586] = 12'h8D0; w_imag[586] = 12'h382;
w_real[587] = 12'h8D6; w_imag[587] = 12'h38D;
w_real[588] = 12'h8DB; w_imag[588] = 12'h398;
w_real[589] = 12'h8E1; w_imag[589] = 12'h3A4;
w_real[590] = 12'h8E7; w_imag[590] = 12'h3AF;
w_real[591] = 12'h8EC; w_imag[591] = 12'h3BA;
w_real[592] = 12'h8F2; w_imag[592] = 12'h3C5;
w_real[593] = 12'h8F8; w_imag[593] = 12'h3D0;
w_real[594] = 12'h8FE; w_imag[594] = 12'h3DB;
w_real[595] = 12'h904; w_imag[595] = 12'h3E6;
w_real[596] = 12'h90B; w_imag[596] = 12'h3F1;
w_real[597] = 12'h911; w_imag[597] = 12'h3FC;
w_real[598] = 12'h917; w_imag[598] = 12'h407;
w_real[599] = 12'h91D; w_imag[599] = 12'h412;
w_real[600] = 12'h924; w_imag[600] = 12'h41C;
w_real[601] = 12'h92A; w_imag[601] = 12'h427;
w_real[602] = 12'h931; w_imag[602] = 12'h432;
w_real[603] = 12'h938; w_imag[603] = 12'h43D;
w_real[604] = 12'h93E; w_imag[604] = 12'h447;
w_real[605] = 12'h945; w_imag[605] = 12'h452;
w_real[606] = 12'h94C; w_imag[606] = 12'h45C;
w_real[607] = 12'h953; w_imag[607] = 12'h467;
w_real[608] = 12'h95A; w_imag[608] = 12'h471;
w_real[609] = 12'h961; w_imag[609] = 12'h47C;
w_real[610] = 12'h968; w_imag[610] = 12'h486;
w_real[611] = 12'h96F; w_imag[611] = 12'h490;
w_real[612] = 12'h976; w_imag[612] = 12'h49B;
w_real[613] = 12'h97D; w_imag[613] = 12'h4A5;
w_real[614] = 12'h985; w_imag[614] = 12'h4AF;
w_real[615] = 12'h98C; w_imag[615] = 12'h4B9;
w_real[616] = 12'h994; w_imag[616] = 12'h4C3;
w_real[617] = 12'h99B; w_imag[617] = 12'h4CE;
w_real[618] = 12'h9A3; w_imag[618] = 12'h4D8;
w_real[619] = 12'h9AA; w_imag[619] = 12'h4E2;
w_real[620] = 12'h9B2; w_imag[620] = 12'h4EB;
w_real[621] = 12'h9BA; w_imag[621] = 12'h4F5;
w_real[622] = 12'h9C2; w_imag[622] = 12'h4FF;
w_real[623] = 12'h9C9; w_imag[623] = 12'h509;
w_real[624] = 12'h9D1; w_imag[624] = 12'h513;
w_real[625] = 12'h9D9; w_imag[625] = 12'h51C;
w_real[626] = 12'h9E1; w_imag[626] = 12'h526;
w_real[627] = 12'h9EA; w_imag[627] = 12'h530;
w_real[628] = 12'h9F2; w_imag[628] = 12'h539;
w_real[629] = 12'h9FA; w_imag[629] = 12'h543;
w_real[630] = 12'hA02; w_imag[630] = 12'h54C;
w_real[631] = 12'hA0B; w_imag[631] = 12'h556;
w_real[632] = 12'hA13; w_imag[632] = 12'h55F;
w_real[633] = 12'hA1B; w_imag[633] = 12'h568;
w_real[634] = 12'hA24; w_imag[634] = 12'h571;
w_real[635] = 12'hA2D; w_imag[635] = 12'h57B;
w_real[636] = 12'hA35; w_imag[636] = 12'h584;
w_real[637] = 12'hA3E; w_imag[637] = 12'h58D;
w_real[638] = 12'hA47; w_imag[638] = 12'h596;
w_real[639] = 12'hA4F; w_imag[639] = 12'h59F;
w_real[640] = 12'hA58; w_imag[640] = 12'h5A8;
w_real[641] = 12'hA61; w_imag[641] = 12'h5B1;
w_real[642] = 12'hA6A; w_imag[642] = 12'h5B9;
w_real[643] = 12'hA73; w_imag[643] = 12'h5C2;
w_real[644] = 12'hA7C; w_imag[644] = 12'h5CB;
w_real[645] = 12'hA85; w_imag[645] = 12'h5D3;
w_real[646] = 12'hA8F; w_imag[646] = 12'h5DC;
w_real[647] = 12'hA98; w_imag[647] = 12'h5E5;
w_real[648] = 12'hAA1; w_imag[648] = 12'h5ED;
w_real[649] = 12'hAAA; w_imag[649] = 12'h5F5;
w_real[650] = 12'hAB4; w_imag[650] = 12'h5FE;
w_real[651] = 12'hABD; w_imag[651] = 12'h606;
w_real[652] = 12'hAC7; w_imag[652] = 12'h60E;
w_real[653] = 12'hAD0; w_imag[653] = 12'h616;
w_real[654] = 12'hADA; w_imag[654] = 12'h61F;
w_real[655] = 12'hAE4; w_imag[655] = 12'h627;
w_real[656] = 12'hAED; w_imag[656] = 12'h62F;
w_real[657] = 12'hAF7; w_imag[657] = 12'h637;
w_real[658] = 12'hB01; w_imag[658] = 12'h63E;
w_real[659] = 12'hB0B; w_imag[659] = 12'h646;
w_real[660] = 12'hB15; w_imag[660] = 12'h64E;
w_real[661] = 12'hB1E; w_imag[661] = 12'h656;
w_real[662] = 12'hB28; w_imag[662] = 12'h65D;
w_real[663] = 12'hB32; w_imag[663] = 12'h665;
w_real[664] = 12'hB3D; w_imag[664] = 12'h66C;
w_real[665] = 12'hB47; w_imag[665] = 12'h674;
w_real[666] = 12'hB51; w_imag[666] = 12'h67B;
w_real[667] = 12'hB5B; w_imag[667] = 12'h683;
w_real[668] = 12'hB65; w_imag[668] = 12'h68A;
w_real[669] = 12'hB70; w_imag[669] = 12'h691;
w_real[670] = 12'hB7A; w_imag[670] = 12'h698;
w_real[671] = 12'hB84; w_imag[671] = 12'h69F;
w_real[672] = 12'hB8F; w_imag[672] = 12'h6A6;
w_real[673] = 12'hB99; w_imag[673] = 12'h6AD;
w_real[674] = 12'hBA4; w_imag[674] = 12'h6B4;
w_real[675] = 12'hBAE; w_imag[675] = 12'h6BB;
w_real[676] = 12'hBB9; w_imag[676] = 12'h6C2;
w_real[677] = 12'hBC3; w_imag[677] = 12'h6C8;
w_real[678] = 12'hBCE; w_imag[678] = 12'h6CF;
w_real[679] = 12'hBD9; w_imag[679] = 12'h6D6;
w_real[680] = 12'hBE4; w_imag[680] = 12'h6DC;
w_real[681] = 12'hBEE; w_imag[681] = 12'h6E3;
w_real[682] = 12'hBF9; w_imag[682] = 12'h6E9;
w_real[683] = 12'hC04; w_imag[683] = 12'h6EF;
w_real[684] = 12'hC0F; w_imag[684] = 12'h6F5;
w_real[685] = 12'hC1A; w_imag[685] = 12'h6FC;
w_real[686] = 12'hC25; w_imag[686] = 12'h702;
w_real[687] = 12'hC30; w_imag[687] = 12'h708;
w_real[688] = 12'hC3B; w_imag[688] = 12'h70E;
w_real[689] = 12'hC46; w_imag[689] = 12'h714;
w_real[690] = 12'hC51; w_imag[690] = 12'h719;
w_real[691] = 12'hC5C; w_imag[691] = 12'h71F;
w_real[692] = 12'hC68; w_imag[692] = 12'h725;
w_real[693] = 12'hC73; w_imag[693] = 12'h72A;
w_real[694] = 12'hC7E; w_imag[694] = 12'h730;
w_real[695] = 12'hC8A; w_imag[695] = 12'h735;
w_real[696] = 12'hC95; w_imag[696] = 12'h73B;
w_real[697] = 12'hCA0; w_imag[697] = 12'h740;
w_real[698] = 12'hCAC; w_imag[698] = 12'h745;
w_real[699] = 12'hCB7; w_imag[699] = 12'h74B;
w_real[700] = 12'hCC3; w_imag[700] = 12'h750;
w_real[701] = 12'hCCE; w_imag[701] = 12'h755;
w_real[702] = 12'hCDA; w_imag[702] = 12'h75A;
w_real[703] = 12'hCE5; w_imag[703] = 12'h75F;
w_real[704] = 12'hCF1; w_imag[704] = 12'h764;
w_real[705] = 12'hCFC; w_imag[705] = 12'h768;
w_real[706] = 12'hD08; w_imag[706] = 12'h76D;
w_real[707] = 12'hD14; w_imag[707] = 12'h772;
w_real[708] = 12'hD1F; w_imag[708] = 12'h776;
w_real[709] = 12'hD2B; w_imag[709] = 12'h77B;
w_real[710] = 12'hD37; w_imag[710] = 12'h77F;
w_real[711] = 12'hD43; w_imag[711] = 12'h784;
w_real[712] = 12'hD4F; w_imag[712] = 12'h788;
w_real[713] = 12'hD5A; w_imag[713] = 12'h78C;
w_real[714] = 12'hD66; w_imag[714] = 12'h790;
w_real[715] = 12'hD72; w_imag[715] = 12'h794;
w_real[716] = 12'hD7E; w_imag[716] = 12'h798;
w_real[717] = 12'hD8A; w_imag[717] = 12'h79C;
w_real[718] = 12'hD96; w_imag[718] = 12'h7A0;
w_real[719] = 12'hDA2; w_imag[719] = 12'h7A4;
w_real[720] = 12'hDAE; w_imag[720] = 12'h7A7;
w_real[721] = 12'hDBA; w_imag[721] = 12'h7AB;
w_real[722] = 12'hDC6; w_imag[722] = 12'h7AE;
w_real[723] = 12'hDD2; w_imag[723] = 12'h7B2;
w_real[724] = 12'hDDE; w_imag[724] = 12'h7B5;
w_real[725] = 12'hDEA; w_imag[725] = 12'h7B9;
w_real[726] = 12'hDF7; w_imag[726] = 12'h7BC;
w_real[727] = 12'hE03; w_imag[727] = 12'h7BF;
w_real[728] = 12'hE0F; w_imag[728] = 12'h7C2;
w_real[729] = 12'hE1B; w_imag[729] = 12'h7C5;
w_real[730] = 12'hE27; w_imag[730] = 12'h7C8;
w_real[731] = 12'hE34; w_imag[731] = 12'h7CB;
w_real[732] = 12'hE40; w_imag[732] = 12'h7CE;
w_real[733] = 12'hE4C; w_imag[733] = 12'h7D0;
w_real[734] = 12'hE58; w_imag[734] = 12'h7D3;
w_real[735] = 12'hE65; w_imag[735] = 12'h7D6;
w_real[736] = 12'hE71; w_imag[736] = 12'h7D8;
w_real[737] = 12'hE7D; w_imag[737] = 12'h7DB;
w_real[738] = 12'hE8A; w_imag[738] = 12'h7DD;
w_real[739] = 12'hE96; w_imag[739] = 12'h7DF;
w_real[740] = 12'hEA2; w_imag[740] = 12'h7E1;
w_real[741] = 12'hEAF; w_imag[741] = 12'h7E3;
w_real[742] = 12'hEBB; w_imag[742] = 12'h7E5;
w_real[743] = 12'hEC8; w_imag[743] = 12'h7E7;
w_real[744] = 12'hED4; w_imag[744] = 12'h7E9;
w_real[745] = 12'hEE0; w_imag[745] = 12'h7EB;
w_real[746] = 12'hEED; w_imag[746] = 12'h7ED;
w_real[747] = 12'hEF9; w_imag[747] = 12'h7EF;
w_real[748] = 12'hF06; w_imag[748] = 12'h7F0;
w_real[749] = 12'hF12; w_imag[749] = 12'h7F2;
w_real[750] = 12'hF1F; w_imag[750] = 12'h7F3;
w_real[751] = 12'hF2B; w_imag[751] = 12'h7F4;
w_real[752] = 12'hF38; w_imag[752] = 12'h7F6;
w_real[753] = 12'hF44; w_imag[753] = 12'h7F7;
w_real[754] = 12'hF51; w_imag[754] = 12'h7F8;
w_real[755] = 12'hF5D; w_imag[755] = 12'h7F9;
w_real[756] = 12'hF6A; w_imag[756] = 12'h7FA;
w_real[757] = 12'hF76; w_imag[757] = 12'h7FB;
w_real[758] = 12'hF83; w_imag[758] = 12'h7FC;
w_real[759] = 12'hF8F; w_imag[759] = 12'h7FC;
w_real[760] = 12'hF9C; w_imag[760] = 12'h7FD;
w_real[761] = 12'hFA9; w_imag[761] = 12'h7FE;
w_real[762] = 12'hFB5; w_imag[762] = 12'h7FE;
w_real[763] = 12'hFC2; w_imag[763] = 12'h7FF;
w_real[764] = 12'hFCE; w_imag[764] = 12'h7FF;
w_real[765] = 12'hFDB; w_imag[765] = 12'h7FF;
w_real[766] = 12'hFE7; w_imag[766] = 12'h7FF;
w_real[767] = 12'hFF4; w_imag[767] = 12'h7FF;
w_real[768] = 12'h000; w_imag[768] = 12'h7FF;
w_real[769] = 12'h00C; w_imag[769] = 12'h7FF;
w_real[770] = 12'h019; w_imag[770] = 12'h7FF;
w_real[771] = 12'h025; w_imag[771] = 12'h7FF;
w_real[772] = 12'h032; w_imag[772] = 12'h7FF;
w_real[773] = 12'h03E; w_imag[773] = 12'h7FF;
w_real[774] = 12'h04B; w_imag[774] = 12'h7FE;
w_real[775] = 12'h057; w_imag[775] = 12'h7FE;
w_real[776] = 12'h064; w_imag[776] = 12'h7FD;
w_real[777] = 12'h071; w_imag[777] = 12'h7FC;
w_real[778] = 12'h07D; w_imag[778] = 12'h7FC;
w_real[779] = 12'h08A; w_imag[779] = 12'h7FB;
w_real[780] = 12'h096; w_imag[780] = 12'h7FA;
w_real[781] = 12'h0A3; w_imag[781] = 12'h7F9;
w_real[782] = 12'h0AF; w_imag[782] = 12'h7F8;
w_real[783] = 12'h0BC; w_imag[783] = 12'h7F7;
w_real[784] = 12'h0C8; w_imag[784] = 12'h7F6;
w_real[785] = 12'h0D5; w_imag[785] = 12'h7F4;
w_real[786] = 12'h0E1; w_imag[786] = 12'h7F3;
w_real[787] = 12'h0EE; w_imag[787] = 12'h7F2;
w_real[788] = 12'h0FA; w_imag[788] = 12'h7F0;
w_real[789] = 12'h107; w_imag[789] = 12'h7EF;
w_real[790] = 12'h113; w_imag[790] = 12'h7ED;
w_real[791] = 12'h120; w_imag[791] = 12'h7EB;
w_real[792] = 12'h12C; w_imag[792] = 12'h7E9;
w_real[793] = 12'h138; w_imag[793] = 12'h7E7;
w_real[794] = 12'h145; w_imag[794] = 12'h7E5;
w_real[795] = 12'h151; w_imag[795] = 12'h7E3;
w_real[796] = 12'h15E; w_imag[796] = 12'h7E1;
w_real[797] = 12'h16A; w_imag[797] = 12'h7DF;
w_real[798] = 12'h176; w_imag[798] = 12'h7DD;
w_real[799] = 12'h183; w_imag[799] = 12'h7DB;
w_real[800] = 12'h18F; w_imag[800] = 12'h7D8;
w_real[801] = 12'h19B; w_imag[801] = 12'h7D6;
w_real[802] = 12'h1A8; w_imag[802] = 12'h7D3;
w_real[803] = 12'h1B4; w_imag[803] = 12'h7D0;
w_real[804] = 12'h1C0; w_imag[804] = 12'h7CE;
w_real[805] = 12'h1CC; w_imag[805] = 12'h7CB;
w_real[806] = 12'h1D9; w_imag[806] = 12'h7C8;
w_real[807] = 12'h1E5; w_imag[807] = 12'h7C5;
w_real[808] = 12'h1F1; w_imag[808] = 12'h7C2;
w_real[809] = 12'h1FD; w_imag[809] = 12'h7BF;
w_real[810] = 12'h209; w_imag[810] = 12'h7BC;
w_real[811] = 12'h216; w_imag[811] = 12'h7B9;
w_real[812] = 12'h222; w_imag[812] = 12'h7B5;
w_real[813] = 12'h22E; w_imag[813] = 12'h7B2;
w_real[814] = 12'h23A; w_imag[814] = 12'h7AE;
w_real[815] = 12'h246; w_imag[815] = 12'h7AB;
w_real[816] = 12'h252; w_imag[816] = 12'h7A7;
w_real[817] = 12'h25E; w_imag[817] = 12'h7A4;
w_real[818] = 12'h26A; w_imag[818] = 12'h7A0;
w_real[819] = 12'h276; w_imag[819] = 12'h79C;
w_real[820] = 12'h282; w_imag[820] = 12'h798;
w_real[821] = 12'h28E; w_imag[821] = 12'h794;
w_real[822] = 12'h29A; w_imag[822] = 12'h790;
w_real[823] = 12'h2A6; w_imag[823] = 12'h78C;
w_real[824] = 12'h2B1; w_imag[824] = 12'h788;
w_real[825] = 12'h2BD; w_imag[825] = 12'h784;
w_real[826] = 12'h2C9; w_imag[826] = 12'h77F;
w_real[827] = 12'h2D5; w_imag[827] = 12'h77B;
w_real[828] = 12'h2E1; w_imag[828] = 12'h776;
w_real[829] = 12'h2EC; w_imag[829] = 12'h772;
w_real[830] = 12'h2F8; w_imag[830] = 12'h76D;
w_real[831] = 12'h304; w_imag[831] = 12'h768;
w_real[832] = 12'h30F; w_imag[832] = 12'h764;
w_real[833] = 12'h31B; w_imag[833] = 12'h75F;
w_real[834] = 12'h326; w_imag[834] = 12'h75A;
w_real[835] = 12'h332; w_imag[835] = 12'h755;
w_real[836] = 12'h33D; w_imag[836] = 12'h750;
w_real[837] = 12'h349; w_imag[837] = 12'h74B;
w_real[838] = 12'h354; w_imag[838] = 12'h745;
w_real[839] = 12'h360; w_imag[839] = 12'h740;
w_real[840] = 12'h36B; w_imag[840] = 12'h73B;
w_real[841] = 12'h376; w_imag[841] = 12'h735;
w_real[842] = 12'h382; w_imag[842] = 12'h730;
w_real[843] = 12'h38D; w_imag[843] = 12'h72A;
w_real[844] = 12'h398; w_imag[844] = 12'h725;
w_real[845] = 12'h3A4; w_imag[845] = 12'h71F;
w_real[846] = 12'h3AF; w_imag[846] = 12'h719;
w_real[847] = 12'h3BA; w_imag[847] = 12'h714;
w_real[848] = 12'h3C5; w_imag[848] = 12'h70E;
w_real[849] = 12'h3D0; w_imag[849] = 12'h708;
w_real[850] = 12'h3DB; w_imag[850] = 12'h702;
w_real[851] = 12'h3E6; w_imag[851] = 12'h6FC;
w_real[852] = 12'h3F1; w_imag[852] = 12'h6F5;
w_real[853] = 12'h3FC; w_imag[853] = 12'h6EF;
w_real[854] = 12'h407; w_imag[854] = 12'h6E9;
w_real[855] = 12'h412; w_imag[855] = 12'h6E3;
w_real[856] = 12'h41C; w_imag[856] = 12'h6DC;
w_real[857] = 12'h427; w_imag[857] = 12'h6D6;
w_real[858] = 12'h432; w_imag[858] = 12'h6CF;
w_real[859] = 12'h43D; w_imag[859] = 12'h6C8;
w_real[860] = 12'h447; w_imag[860] = 12'h6C2;
w_real[861] = 12'h452; w_imag[861] = 12'h6BB;
w_real[862] = 12'h45C; w_imag[862] = 12'h6B4;
w_real[863] = 12'h467; w_imag[863] = 12'h6AD;
w_real[864] = 12'h471; w_imag[864] = 12'h6A6;
w_real[865] = 12'h47C; w_imag[865] = 12'h69F;
w_real[866] = 12'h486; w_imag[866] = 12'h698;
w_real[867] = 12'h490; w_imag[867] = 12'h691;
w_real[868] = 12'h49B; w_imag[868] = 12'h68A;
w_real[869] = 12'h4A5; w_imag[869] = 12'h683;
w_real[870] = 12'h4AF; w_imag[870] = 12'h67B;
w_real[871] = 12'h4B9; w_imag[871] = 12'h674;
w_real[872] = 12'h4C3; w_imag[872] = 12'h66C;
w_real[873] = 12'h4CE; w_imag[873] = 12'h665;
w_real[874] = 12'h4D8; w_imag[874] = 12'h65D;
w_real[875] = 12'h4E2; w_imag[875] = 12'h656;
w_real[876] = 12'h4EB; w_imag[876] = 12'h64E;
w_real[877] = 12'h4F5; w_imag[877] = 12'h646;
w_real[878] = 12'h4FF; w_imag[878] = 12'h63E;
w_real[879] = 12'h509; w_imag[879] = 12'h637;
w_real[880] = 12'h513; w_imag[880] = 12'h62F;
w_real[881] = 12'h51C; w_imag[881] = 12'h627;
w_real[882] = 12'h526; w_imag[882] = 12'h61F;
w_real[883] = 12'h530; w_imag[883] = 12'h616;
w_real[884] = 12'h539; w_imag[884] = 12'h60E;
w_real[885] = 12'h543; w_imag[885] = 12'h606;
w_real[886] = 12'h54C; w_imag[886] = 12'h5FE;
w_real[887] = 12'h556; w_imag[887] = 12'h5F5;
w_real[888] = 12'h55F; w_imag[888] = 12'h5ED;
w_real[889] = 12'h568; w_imag[889] = 12'h5E5;
w_real[890] = 12'h571; w_imag[890] = 12'h5DC;
w_real[891] = 12'h57B; w_imag[891] = 12'h5D3;
w_real[892] = 12'h584; w_imag[892] = 12'h5CB;
w_real[893] = 12'h58D; w_imag[893] = 12'h5C2;
w_real[894] = 12'h596; w_imag[894] = 12'h5B9;
w_real[895] = 12'h59F; w_imag[895] = 12'h5B1;
w_real[896] = 12'h5A8; w_imag[896] = 12'h5A8;
w_real[897] = 12'h5B1; w_imag[897] = 12'h59F;
w_real[898] = 12'h5B9; w_imag[898] = 12'h596;
w_real[899] = 12'h5C2; w_imag[899] = 12'h58D;
w_real[900] = 12'h5CB; w_imag[900] = 12'h584;
w_real[901] = 12'h5D3; w_imag[901] = 12'h57B;
w_real[902] = 12'h5DC; w_imag[902] = 12'h571;
w_real[903] = 12'h5E5; w_imag[903] = 12'h568;
w_real[904] = 12'h5ED; w_imag[904] = 12'h55F;
w_real[905] = 12'h5F5; w_imag[905] = 12'h556;
w_real[906] = 12'h5FE; w_imag[906] = 12'h54C;
w_real[907] = 12'h606; w_imag[907] = 12'h543;
w_real[908] = 12'h60E; w_imag[908] = 12'h539;
w_real[909] = 12'h616; w_imag[909] = 12'h530;
w_real[910] = 12'h61F; w_imag[910] = 12'h526;
w_real[911] = 12'h627; w_imag[911] = 12'h51C;
w_real[912] = 12'h62F; w_imag[912] = 12'h513;
w_real[913] = 12'h637; w_imag[913] = 12'h509;
w_real[914] = 12'h63E; w_imag[914] = 12'h4FF;
w_real[915] = 12'h646; w_imag[915] = 12'h4F5;
w_real[916] = 12'h64E; w_imag[916] = 12'h4EB;
w_real[917] = 12'h656; w_imag[917] = 12'h4E2;
w_real[918] = 12'h65D; w_imag[918] = 12'h4D8;
w_real[919] = 12'h665; w_imag[919] = 12'h4CE;
w_real[920] = 12'h66C; w_imag[920] = 12'h4C3;
w_real[921] = 12'h674; w_imag[921] = 12'h4B9;
w_real[922] = 12'h67B; w_imag[922] = 12'h4AF;
w_real[923] = 12'h683; w_imag[923] = 12'h4A5;
w_real[924] = 12'h68A; w_imag[924] = 12'h49B;
w_real[925] = 12'h691; w_imag[925] = 12'h490;
w_real[926] = 12'h698; w_imag[926] = 12'h486;
w_real[927] = 12'h69F; w_imag[927] = 12'h47C;
w_real[928] = 12'h6A6; w_imag[928] = 12'h471;
w_real[929] = 12'h6AD; w_imag[929] = 12'h467;
w_real[930] = 12'h6B4; w_imag[930] = 12'h45C;
w_real[931] = 12'h6BB; w_imag[931] = 12'h452;
w_real[932] = 12'h6C2; w_imag[932] = 12'h447;
w_real[933] = 12'h6C8; w_imag[933] = 12'h43D;
w_real[934] = 12'h6CF; w_imag[934] = 12'h432;
w_real[935] = 12'h6D6; w_imag[935] = 12'h427;
w_real[936] = 12'h6DC; w_imag[936] = 12'h41C;
w_real[937] = 12'h6E3; w_imag[937] = 12'h412;
w_real[938] = 12'h6E9; w_imag[938] = 12'h407;
w_real[939] = 12'h6EF; w_imag[939] = 12'h3FC;
w_real[940] = 12'h6F5; w_imag[940] = 12'h3F1;
w_real[941] = 12'h6FC; w_imag[941] = 12'h3E6;
w_real[942] = 12'h702; w_imag[942] = 12'h3DB;
w_real[943] = 12'h708; w_imag[943] = 12'h3D0;
w_real[944] = 12'h70E; w_imag[944] = 12'h3C5;
w_real[945] = 12'h714; w_imag[945] = 12'h3BA;
w_real[946] = 12'h719; w_imag[946] = 12'h3AF;
w_real[947] = 12'h71F; w_imag[947] = 12'h3A4;
w_real[948] = 12'h725; w_imag[948] = 12'h398;
w_real[949] = 12'h72A; w_imag[949] = 12'h38D;
w_real[950] = 12'h730; w_imag[950] = 12'h382;
w_real[951] = 12'h735; w_imag[951] = 12'h376;
w_real[952] = 12'h73B; w_imag[952] = 12'h36B;
w_real[953] = 12'h740; w_imag[953] = 12'h360;
w_real[954] = 12'h745; w_imag[954] = 12'h354;
w_real[955] = 12'h74B; w_imag[955] = 12'h349;
w_real[956] = 12'h750; w_imag[956] = 12'h33D;
w_real[957] = 12'h755; w_imag[957] = 12'h332;
w_real[958] = 12'h75A; w_imag[958] = 12'h326;
w_real[959] = 12'h75F; w_imag[959] = 12'h31B;
w_real[960] = 12'h764; w_imag[960] = 12'h30F;
w_real[961] = 12'h768; w_imag[961] = 12'h304;
w_real[962] = 12'h76D; w_imag[962] = 12'h2F8;
w_real[963] = 12'h772; w_imag[963] = 12'h2EC;
w_real[964] = 12'h776; w_imag[964] = 12'h2E1;
w_real[965] = 12'h77B; w_imag[965] = 12'h2D5;
w_real[966] = 12'h77F; w_imag[966] = 12'h2C9;
w_real[967] = 12'h784; w_imag[967] = 12'h2BD;
w_real[968] = 12'h788; w_imag[968] = 12'h2B1;
w_real[969] = 12'h78C; w_imag[969] = 12'h2A6;
w_real[970] = 12'h790; w_imag[970] = 12'h29A;
w_real[971] = 12'h794; w_imag[971] = 12'h28E;
w_real[972] = 12'h798; w_imag[972] = 12'h282;
w_real[973] = 12'h79C; w_imag[973] = 12'h276;
w_real[974] = 12'h7A0; w_imag[974] = 12'h26A;
w_real[975] = 12'h7A4; w_imag[975] = 12'h25E;
w_real[976] = 12'h7A7; w_imag[976] = 12'h252;
w_real[977] = 12'h7AB; w_imag[977] = 12'h246;
w_real[978] = 12'h7AE; w_imag[978] = 12'h23A;
w_real[979] = 12'h7B2; w_imag[979] = 12'h22E;
w_real[980] = 12'h7B5; w_imag[980] = 12'h222;
w_real[981] = 12'h7B9; w_imag[981] = 12'h216;
w_real[982] = 12'h7BC; w_imag[982] = 12'h209;
w_real[983] = 12'h7BF; w_imag[983] = 12'h1FD;
w_real[984] = 12'h7C2; w_imag[984] = 12'h1F1;
w_real[985] = 12'h7C5; w_imag[985] = 12'h1E5;
w_real[986] = 12'h7C8; w_imag[986] = 12'h1D9;
w_real[987] = 12'h7CB; w_imag[987] = 12'h1CC;
w_real[988] = 12'h7CE; w_imag[988] = 12'h1C0;
w_real[989] = 12'h7D0; w_imag[989] = 12'h1B4;
w_real[990] = 12'h7D3; w_imag[990] = 12'h1A8;
w_real[991] = 12'h7D6; w_imag[991] = 12'h19B;
w_real[992] = 12'h7D8; w_imag[992] = 12'h18F;
w_real[993] = 12'h7DB; w_imag[993] = 12'h183;
w_real[994] = 12'h7DD; w_imag[994] = 12'h176;
w_real[995] = 12'h7DF; w_imag[995] = 12'h16A;
w_real[996] = 12'h7E1; w_imag[996] = 12'h15E;
w_real[997] = 12'h7E3; w_imag[997] = 12'h151;
w_real[998] = 12'h7E5; w_imag[998] = 12'h145;
w_real[999] = 12'h7E7; w_imag[999] = 12'h138;
w_real[1000] = 12'h7E9; w_imag[1000] = 12'h12C;
w_real[1001] = 12'h7EB; w_imag[1001] = 12'h120;
w_real[1002] = 12'h7ED; w_imag[1002] = 12'h113;
w_real[1003] = 12'h7EF; w_imag[1003] = 12'h107;
w_real[1004] = 12'h7F0; w_imag[1004] = 12'h0FA;
w_real[1005] = 12'h7F2; w_imag[1005] = 12'h0EE;
w_real[1006] = 12'h7F3; w_imag[1006] = 12'h0E1;
w_real[1007] = 12'h7F4; w_imag[1007] = 12'h0D5;
w_real[1008] = 12'h7F6; w_imag[1008] = 12'h0C8;
w_real[1009] = 12'h7F7; w_imag[1009] = 12'h0BC;
w_real[1010] = 12'h7F8; w_imag[1010] = 12'h0AF;
w_real[1011] = 12'h7F9; w_imag[1011] = 12'h0A3;
w_real[1012] = 12'h7FA; w_imag[1012] = 12'h096;
w_real[1013] = 12'h7FB; w_imag[1013] = 12'h08A;
w_real[1014] = 12'h7FC; w_imag[1014] = 12'h07D;
w_real[1015] = 12'h7FC; w_imag[1015] = 12'h071;
w_real[1016] = 12'h7FD; w_imag[1016] = 12'h064;
w_real[1017] = 12'h7FE; w_imag[1017] = 12'h057;
w_real[1018] = 12'h7FE; w_imag[1018] = 12'h04B;
w_real[1019] = 12'h7FF; w_imag[1019] = 12'h03E;
w_real[1020] = 12'h7FF; w_imag[1020] = 12'h032;
w_real[1021] = 12'h7FF; w_imag[1021] = 12'h025;
w_real[1022] = 12'h7FF; w_imag[1022] = 12'h019;
w_real[1023] = 12'h7FF; w_imag[1023] = 12'h00C;
