gen_input_real[0] = 24'sd0;
gen_input_real[16] = 24'sd2047;
gen_input_real[32] = -24'sd420;
gen_input_real[48] = -24'sd1519;
gen_input_real[4] = 24'sd609;
gen_input_real[20] = 24'sd950;
gen_input_real[36] = -24'sd628;
gen_input_real[52] = -24'sd494;
gen_input_real[8] = 24'sd669;
gen_input_real[24] = 24'sd223;
gen_input_real[40] = -24'sd736;
gen_input_real[56] = -24'sd120;
gen_input_real[12] = 24'sd681;
gen_input_real[28] = 24'sd59;
gen_input_real[44] = -24'sd454;
gen_input_real[60] = -24'sd89;
gen_input_real[1] = 24'sd137;
gen_input_real[17] = 24'sd159;
gen_input_real[33] = 24'sd150;
gen_input_real[49] = -24'sd120;
gen_input_real[5] = -24'sd277;
gen_input_real[21] = -24'sd43;
gen_input_real[37] = 24'sd258;
gen_input_real[53] = 24'sd268;
gen_input_real[9] = -24'sd236;
gen_input_real[25] = -24'sd406;
gen_input_real[41] = 24'sd217;
gen_input_real[57] = 24'sd282;
gen_input_real[13] = -24'sd133;
gen_input_real[29] = 24'sd37;
gen_input_real[45] = -24'sd48;
gen_input_real[61] = -24'sd189;
gen_input_real[2] = 24'sd189;
gen_input_real[18] = 24'sd48;
gen_input_real[34] = -24'sd37;
gen_input_real[50] = 24'sd133;
gen_input_real[6] = -24'sd282;
gen_input_real[22] = -24'sd217;
gen_input_real[38] = 24'sd406;
gen_input_real[54] = 24'sd236;
gen_input_real[10] = -24'sd268;
gen_input_real[26] = -24'sd258;
gen_input_real[42] = 24'sd43;
gen_input_real[58] = 24'sd277;
gen_input_real[14] = 24'sd120;
gen_input_real[30] = -24'sd150;
gen_input_real[46] = -24'sd159;
gen_input_real[62] = -24'sd137;
gen_input_real[3] = 24'sd89;
gen_input_real[19] = 24'sd454;
gen_input_real[35] = -24'sd59;
gen_input_real[51] = -24'sd681;
gen_input_real[7] = 24'sd120;
gen_input_real[23] = 24'sd736;
gen_input_real[39] = -24'sd223;
gen_input_real[55] = -24'sd669;
gen_input_real[11] = 24'sd494;
gen_input_real[27] = 24'sd628;
gen_input_real[43] = -24'sd950;
gen_input_real[59] = -24'sd609;
gen_input_real[15] = 24'sd1519;
gen_input_real[31] = 24'sd420;
gen_input_real[47] = -24'sd2047;
gen_input_real[63] = 24'sd0;
