0 0
0 -6
0 -4
0 -3
0 -6
0 -10
0 -10
1 -12
1 -10
2 -25
1 -15
2 -21
5 -34
1 -12
4 -25
4 -24
8 -44
6 -32
7 -35
10 -42
18 -73
8 -30
13 -50
15 -54
32 -108
12 -39
17 -53
21 -62
26 -73
30 -82
30 -79
33 -84
30 -73
41 -96
58 -131
68 -149
301 -636
8 -16
36 -71
60 -116
82 -155
308 -560
45 -79
338 -580
-19 33
26 -42
45 -72
73 -112
86 -128
117 -171
136 -193
209 -289
852 -1149
-69 91
60 -77
119 -149
172 -209
243 -289
335 -388
552 -624
1953 -2155
1455 -1566
1010 -1061
-873 894
-447 447
-291 284
-209 199
-141 131
-81 73
-26 23
47 -40
155 -131
394 -323
2178 -1743
-999 779
-448 341
-272 201
-108 78
552 -389
-571 391
-344 230
-258 168
-227 144
-195 120
-143 85
-89 51
234 -132
-367 202
-212 113
-142 73
84 -42
-333 162
-231 109
-176 80
-128 56
1 0
-214 88
42 -16
-350 135
-244 90
-227 81
-191 65
-175 58
-128 40
-219 66
-184 53
-173 48
-167 44
-150 37
-182 43
-158 35
-158 33
-174 34
-149 27
-156 27
-155 24
-155 23
-148 20
-157 19
-151 16
-147 14
-143 12
-153 11
-144 8
-147 7
-147 5
-152 3
-146 1
-146 0
-146 -1
-152 -3
-147 -5
-147 -7
-144 -8
-153 -11
-143 -12
-147 -14
-151 -16
-157 -19
-148 -20
-155 -23
-155 -24
-156 -27
-149 -27
-174 -34
-158 -33
-158 -35
-182 -43
-150 -37
-167 -44
-173 -48
-184 -53
-219 -66
-128 -40
-175 -58
-191 -65
-227 -81
-244 -90
-350 -135
42 16
-214 -88
1 0
-128 -56
-176 -80
-231 -109
-333 -162
84 42
-142 -73
-212 -113
-367 -202
234 132
-89 -51
-143 -85
-195 -120
-227 -144
-258 -168
-344 -230
-571 -391
552 389
-108 -78
-272 -201
-448 -341
-999 -779
2178 1743
394 323
155 131
47 40
-26 -23
-81 -73
-141 -131
-209 -199
-291 -284
-447 -447
-873 -894
1010 1061
1455 1566
1953 2155
552 624
335 388
243 289
172 209
119 149
60 77
-69 -91
852 1149
209 289
136 193
117 171
86 128
73 112
45 72
26 42
-19 -33
338 580
45 79
308 560
82 155
60 116
36 71
8 16
301 636
68 149
58 131
41 96
30 73
33 84
30 79
30 82
26 73
21 62
17 53
12 39
32 108
15 54
13 50
8 30
18 73
10 42
7 35
6 32
8 44
4 24
4 25
1 12
5 34
2 21
1 15
2 25
1 10
1 12
0 10
0 10
0 6
0 3
0 4
0 6
