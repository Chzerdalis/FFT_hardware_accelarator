0 0
0 -29
1 -53
3 -86
5 -109
9 -148
12 -163
18 -216
22 -224
28 -259
39 -320
44 -324
63 -429
61 -379
73 -422
87 -468
136 -686
108 -510
126 -561
150 -632
277 -1106
174 -662
199 -721
237 -819
523 -1726
235 -743
282 -855
321 -934
358 -1001
411 -1106
457 -1185
520 -1300
582 -1405
683 -1594
830 -1872
1137 -2484
4885 -10329
105 -216
603 -1198
906 -1747
1337 -2503
4949 -8992
689 -1216
5444 -9341
-270 452
464 -753
807 -1274
1106 -1701
1404 -2102
1768 -2577
2300 -3267
3465 -4794
13871 -18703
-1202 1580
909 -1165
1874 -2341
2752 -3353
3847 -4573
5519 -6398
9030 -10212
31642 -34912
23749 -25565
16505 -17336
-14301 14656
-7262 7262
-4765 4649
-3339 3179
-2309 2145
-1417 1284
-510 451
614 -530
2364 -1989
6297 -5168
35688 -28563
-16423 12817
-7258 5522
-4304 3192
-1776 1284
8995 -6335
-9385 6439
-5570 3721
-4335 2820
-3601 2280
-3016 1858
-2372 1422
-1364 795
3913 -2217
-5906 3251
-3493 1867
-2335 1211
1389 -699
-5328 2600
-3557 1682
-2867 1313
-2191 971
61 -26
-3448 1428
513 -205
-5642 2176
-3927 1459
-3425 1225
-3121 1073
-2851 942
-2121 672
-3439 1043
-2972 862
-2822 781
-2678 705
-2365 592
-2898 688
-2666 598
-2472 523
-2743 545
-2595 483
-2555 443
-2474 398
-2541 376
-2488 337
-2468 304
-2435 270
-2433 239
-2421 208
-2412 177
-2390 146
-2386 117
-2381 87
-2383 58
-2377 29
-2392 0
-2377 -29
-2383 -58
-2381 -87
-2386 -117
-2390 -146
-2412 -177
-2421 -208
-2433 -239
-2435 -270
-2468 -304
-2488 -337
-2541 -376
-2474 -398
-2555 -443
-2595 -483
-2743 -545
-2472 -523
-2666 -598
-2898 -688
-2365 -592
-2678 -705
-2822 -781
-2972 -862
-3439 -1043
-2121 -672
-2851 -942
-3121 -1073
-3425 -1225
-3927 -1459
-5642 -2176
513 205
-3448 -1428
61 26
-2191 -971
-2867 -1313
-3557 -1682
-5328 -2600
1389 699
-2335 -1211
-3493 -1867
-5906 -3251
3913 2217
-1364 -795
-2372 -1422
-3016 -1858
-3601 -2280
-4335 -2820
-5570 -3721
-9385 -6439
8995 6335
-1776 -1284
-4304 -3192
-7258 -5522
-16423 -12817
35688 28563
6297 5168
2364 1989
614 530
-510 -451
-1417 -1284
-2309 -2145
-3339 -3179
-4765 -4649
-7262 -7262
-14301 -14656
16505 17336
23749 25565
31642 34912
9030 10212
5519 6398
3847 4573
2752 3353
1874 2341
909 1165
-1202 -1580
13871 18703
3465 4794
2300 3267
1768 2577
1404 2102
1106 1701
807 1274
464 753
-270 -452
5444 9341
689 1216
4949 8992
1337 2503
906 1747
603 1198
105 216
4885 10329
1137 2484
830 1872
683 1594
582 1405
520 1300
457 1185
411 1106
358 1001
321 934
282 855
235 743
523 1726
237 819
199 721
174 662
277 1106
150 632
126 561
108 510
136 686
87 468
73 422
61 379
63 429
44 324
39 320
28 259
22 224
18 216
12 163
9 148
5 109
3 86
1 53
0 29
