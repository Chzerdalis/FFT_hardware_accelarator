0 0
0 2
0 4
0 -15
0 -17
0 -14
0 -6
1 -14
1 -12
2 -18
2 -20
2 -20
3 -21
4 -24
6 -34
4 -26
6 -30
8 -38
9 -42
8 -34
9 -39
12 -48
16 -59
12 -43
13 -43
15 -48
17 -54
21 -62
21 -59
24 -65
30 -79
63 -159
30 -73
36 -85
45 -101
115 -251
109 -232
105 -216
17 -34
35 -69
41 -78
48 -88
54 -96
64 -111
81 -135
87 -142
99 -156
120 -185
142 -213
195 -285
546 -775
463 -641
401 -540
-53 70
55 -71
97 -121
154 -188
223 -265
354 -410
1055 -1193
763 -842
-133 144
119 -125
302 -309
595 -595
2454 -2395
633 -602
1233 -1146
-915 829
254 -224
-734 633
-447 376
-341 280
-263 210
-160 125
-35 26
792 -587
-681 492
-404 284
-324 222
-278 186
-251 163
-228 144
-200 123
-196 117
-182 106
-147 83
-122 67
34 -18
-228 118
-39 19
-256 125
-91 43
-260 119
-223 99
-195 83
-180 74
-176 70
-176 67
-164 61
-126 45
-196 67
-173 57
-161 51
-152 46
-154 44
-150 41
-154 40
-150 37
-154 36
-136 30
-138 29
-142 28
-140 26
-159 27
-150 24
-150 22
-139 18
-149 18
-135 15
-142 14
-139 12
-140 10
-137 8
-136 6
-130 4
-137 3
-140 1
-138 0
-140 -1
-137 -3
-130 -4
-136 -6
-137 -8
-140 -10
-139 -12
-142 -14
-135 -15
-149 -18
-139 -18
-150 -22
-150 -24
-159 -27
-140 -26
-142 -28
-138 -29
-136 -30
-154 -36
-150 -37
-154 -40
-150 -41
-154 -44
-152 -46
-161 -51
-173 -57
-196 -67
-126 -45
-164 -61
-176 -67
-176 -70
-180 -74
-195 -83
-223 -99
-260 -119
-91 -43
-256 -125
-39 -19
-228 -118
34 18
-122 -67
-147 -83
-182 -106
-196 -117
-200 -123
-228 -144
-251 -163
-278 -186
-324 -222
-404 -284
-681 -492
792 587
-35 -26
-160 -125
-263 -210
-341 -280
-447 -376
-734 -633
254 224
-915 -829
1233 1146
633 602
2454 2395
595 595
302 309
119 125
-133 -144
763 842
1055 1193
354 410
223 265
154 188
97 121
55 71
-53 -70
401 540
463 641
546 775
195 285
142 213
120 185
99 156
87 142
81 135
64 111
54 96
48 88
41 78
35 69
17 34
105 216
109 232
115 251
45 101
36 85
30 73
63 159
30 79
24 65
21 59
21 62
17 54
15 48
13 43
12 43
16 59
12 48
9 39
8 34
9 42
8 38
6 30
4 26
6 34
4 24
3 21
2 20
2 20
2 18
1 12
1 14
0 6
0 14
0 17
0 15
0 -4
0 -2
