0 0
0 -4
1 -10
3 -20
6 -31
10 -41
22 -75
20 -58
30 -74
48 -102
75 -141
229 -383
349 -523
56 -76
489 -595
259 -286
329 -329
399 -362
-152 125
-320 237
-211 141
-159 95
-74 39
-86 40
-162 67
-208 74
-163 49
-146 36
-148 29
-145 21
-142 14
-137 6
-146 0
-137 -6
-142 -14
-145 -21
-148 -29
-146 -36
-163 -49
-208 -74
-162 -67
-86 -40
-74 -39
-159 -95
-211 -141
-320 -237
-152 -125
399 362
329 329
259 286
489 595
56 76
349 523
229 383
75 141
48 102
30 74
20 58
22 75
10 41
6 31
3 20
1 10
0 4
