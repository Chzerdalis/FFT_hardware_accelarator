w_real[0] = 16'h7FFF; w_imag[0] = 16'h0000;
w_real[1] = 16'h7FF6; w_imag[1] = 16'hFCDC;
w_real[2] = 16'h7FD8; w_imag[2] = 16'hF9B9;
w_real[3] = 16'h7FA7; w_imag[3] = 16'hF696;
w_real[4] = 16'h7F62; w_imag[4] = 16'hF375;
w_real[5] = 16'h7F09; w_imag[5] = 16'hF055;
w_real[6] = 16'h7E9D; w_imag[6] = 16'hED38;
w_real[7] = 16'h7E1D; w_imag[7] = 16'hEA1E;
w_real[8] = 16'h7D8A; w_imag[8] = 16'hE708;
w_real[9] = 16'h7CE3; w_imag[9] = 16'hE3F5;
w_real[10] = 16'h7C29; w_imag[10] = 16'hE0E7;
w_real[11] = 16'h7B5D; w_imag[11] = 16'hDDDD;
w_real[12] = 16'h7A7D; w_imag[12] = 16'hDAD8;
w_real[13] = 16'h798A; w_imag[13] = 16'hD7DA;
w_real[14] = 16'h7884; w_imag[14] = 16'hD4E1;
w_real[15] = 16'h776C; w_imag[15] = 16'hD1EF;
w_real[16] = 16'h7641; w_imag[16] = 16'hCF05;
w_real[17] = 16'h7504; w_imag[17] = 16'hCC22;
w_real[18] = 16'h73B5; w_imag[18] = 16'hC946;
w_real[19] = 16'h7255; w_imag[19] = 16'hC674;
w_real[20] = 16'h70E2; w_imag[20] = 16'hC3AA;
w_real[21] = 16'h6F5F; w_imag[21] = 16'hC0E9;
w_real[22] = 16'h6DCA; w_imag[22] = 16'hBE32;
w_real[23] = 16'h6C24; w_imag[23] = 16'hBB86;
w_real[24] = 16'h6A6D; w_imag[24] = 16'hB8E4;
w_real[25] = 16'h68A6; w_imag[25] = 16'hB64C;
w_real[26] = 16'h66CF; w_imag[26] = 16'hB3C1;
w_real[27] = 16'h64E8; w_imag[27] = 16'hB141;
w_real[28] = 16'h62F2; w_imag[28] = 16'hAECD;
w_real[29] = 16'h60EC; w_imag[29] = 16'hAC65;
w_real[30] = 16'h5ED7; w_imag[30] = 16'hAA0B;
w_real[31] = 16'h5CB4; w_imag[31] = 16'hA7BE;
w_real[32] = 16'h5A82; w_imag[32] = 16'hA57E;
w_real[33] = 16'h5842; w_imag[33] = 16'hA34C;
w_real[34] = 16'h55F5; w_imag[34] = 16'hA129;
w_real[35] = 16'h539B; w_imag[35] = 16'h9F14;
w_real[36] = 16'h5133; w_imag[36] = 16'h9D0E;
w_real[37] = 16'h4EBF; w_imag[37] = 16'h9B18;
w_real[38] = 16'h4C3F; w_imag[38] = 16'h9931;
w_real[39] = 16'h49B4; w_imag[39] = 16'h975A;
w_real[40] = 16'h471C; w_imag[40] = 16'h9593;
w_real[41] = 16'h447A; w_imag[41] = 16'h93DC;
w_real[42] = 16'h41CE; w_imag[42] = 16'h9236;
w_real[43] = 16'h3F17; w_imag[43] = 16'h90A1;
w_real[44] = 16'h3C56; w_imag[44] = 16'h8F1E;
w_real[45] = 16'h398C; w_imag[45] = 16'h8DAB;
w_real[46] = 16'h36BA; w_imag[46] = 16'h8C4B;
w_real[47] = 16'h33DE; w_imag[47] = 16'h8AFC;
w_real[48] = 16'h30FB; w_imag[48] = 16'h89BF;
w_real[49] = 16'h2E11; w_imag[49] = 16'h8894;
w_real[50] = 16'h2B1F; w_imag[50] = 16'h877C;
w_real[51] = 16'h2826; w_imag[51] = 16'h8676;
w_real[52] = 16'h2528; w_imag[52] = 16'h8583;
w_real[53] = 16'h2223; w_imag[53] = 16'h84A3;
w_real[54] = 16'h1F19; w_imag[54] = 16'h83D7;
w_real[55] = 16'h1C0B; w_imag[55] = 16'h831D;
w_real[56] = 16'h18F8; w_imag[56] = 16'h8276;
w_real[57] = 16'h15E2; w_imag[57] = 16'h81E3;
w_real[58] = 16'h12C8; w_imag[58] = 16'h8163;
w_real[59] = 16'h0FAB; w_imag[59] = 16'h80F7;
w_real[60] = 16'h0C8B; w_imag[60] = 16'h809E;
w_real[61] = 16'h096A; w_imag[61] = 16'h8059;
w_real[62] = 16'h0647; w_imag[62] = 16'h8028;
w_real[63] = 16'h0324; w_imag[63] = 16'h800A;
w_real[64] = 16'h0000; w_imag[64] = 16'h8000;
w_real[65] = 16'hFCDC; w_imag[65] = 16'h800A;
w_real[66] = 16'hF9B9; w_imag[66] = 16'h8028;
w_real[67] = 16'hF696; w_imag[67] = 16'h8059;
w_real[68] = 16'hF375; w_imag[68] = 16'h809E;
w_real[69] = 16'hF055; w_imag[69] = 16'h80F7;
w_real[70] = 16'hED38; w_imag[70] = 16'h8163;
w_real[71] = 16'hEA1E; w_imag[71] = 16'h81E3;
w_real[72] = 16'hE708; w_imag[72] = 16'h8276;
w_real[73] = 16'hE3F5; w_imag[73] = 16'h831D;
w_real[74] = 16'hE0E7; w_imag[74] = 16'h83D7;
w_real[75] = 16'hDDDD; w_imag[75] = 16'h84A3;
w_real[76] = 16'hDAD8; w_imag[76] = 16'h8583;
w_real[77] = 16'hD7DA; w_imag[77] = 16'h8676;
w_real[78] = 16'hD4E1; w_imag[78] = 16'h877C;
w_real[79] = 16'hD1EF; w_imag[79] = 16'h8894;
w_real[80] = 16'hCF05; w_imag[80] = 16'h89BF;
w_real[81] = 16'hCC22; w_imag[81] = 16'h8AFC;
w_real[82] = 16'hC946; w_imag[82] = 16'h8C4B;
w_real[83] = 16'hC674; w_imag[83] = 16'h8DAB;
w_real[84] = 16'hC3AA; w_imag[84] = 16'h8F1E;
w_real[85] = 16'hC0E9; w_imag[85] = 16'h90A1;
w_real[86] = 16'hBE32; w_imag[86] = 16'h9236;
w_real[87] = 16'hBB86; w_imag[87] = 16'h93DC;
w_real[88] = 16'hB8E4; w_imag[88] = 16'h9593;
w_real[89] = 16'hB64C; w_imag[89] = 16'h975A;
w_real[90] = 16'hB3C1; w_imag[90] = 16'h9931;
w_real[91] = 16'hB141; w_imag[91] = 16'h9B18;
w_real[92] = 16'hAECD; w_imag[92] = 16'h9D0E;
w_real[93] = 16'hAC65; w_imag[93] = 16'h9F14;
w_real[94] = 16'hAA0B; w_imag[94] = 16'hA129;
w_real[95] = 16'hA7BE; w_imag[95] = 16'hA34C;
w_real[96] = 16'hA57E; w_imag[96] = 16'hA57E;
w_real[97] = 16'hA34C; w_imag[97] = 16'hA7BE;
w_real[98] = 16'hA129; w_imag[98] = 16'hAA0B;
w_real[99] = 16'h9F14; w_imag[99] = 16'hAC65;
w_real[100] = 16'h9D0E; w_imag[100] = 16'hAECD;
w_real[101] = 16'h9B18; w_imag[101] = 16'hB141;
w_real[102] = 16'h9931; w_imag[102] = 16'hB3C1;
w_real[103] = 16'h975A; w_imag[103] = 16'hB64C;
w_real[104] = 16'h9593; w_imag[104] = 16'hB8E4;
w_real[105] = 16'h93DC; w_imag[105] = 16'hBB86;
w_real[106] = 16'h9236; w_imag[106] = 16'hBE32;
w_real[107] = 16'h90A1; w_imag[107] = 16'hC0E9;
w_real[108] = 16'h8F1E; w_imag[108] = 16'hC3AA;
w_real[109] = 16'h8DAB; w_imag[109] = 16'hC674;
w_real[110] = 16'h8C4B; w_imag[110] = 16'hC946;
w_real[111] = 16'h8AFC; w_imag[111] = 16'hCC22;
w_real[112] = 16'h89BF; w_imag[112] = 16'hCF05;
w_real[113] = 16'h8894; w_imag[113] = 16'hD1EF;
w_real[114] = 16'h877C; w_imag[114] = 16'hD4E1;
w_real[115] = 16'h8676; w_imag[115] = 16'hD7DA;
w_real[116] = 16'h8583; w_imag[116] = 16'hDAD8;
w_real[117] = 16'h84A3; w_imag[117] = 16'hDDDD;
w_real[118] = 16'h83D7; w_imag[118] = 16'hE0E7;
w_real[119] = 16'h831D; w_imag[119] = 16'hE3F5;
w_real[120] = 16'h8276; w_imag[120] = 16'hE708;
w_real[121] = 16'h81E3; w_imag[121] = 16'hEA1E;
w_real[122] = 16'h8163; w_imag[122] = 16'hED38;
w_real[123] = 16'h80F7; w_imag[123] = 16'hF055;
w_real[124] = 16'h809E; w_imag[124] = 16'hF375;
w_real[125] = 16'h8059; w_imag[125] = 16'hF696;
w_real[126] = 16'h8028; w_imag[126] = 16'hF9B9;
w_real[127] = 16'h800A; w_imag[127] = 16'hFCDC;
w_real[128] = 16'h8000; w_imag[128] = 16'h0000;
w_real[129] = 16'h800A; w_imag[129] = 16'h0324;
w_real[130] = 16'h8028; w_imag[130] = 16'h0647;
w_real[131] = 16'h8059; w_imag[131] = 16'h096A;
w_real[132] = 16'h809E; w_imag[132] = 16'h0C8B;
w_real[133] = 16'h80F7; w_imag[133] = 16'h0FAB;
w_real[134] = 16'h8163; w_imag[134] = 16'h12C8;
w_real[135] = 16'h81E3; w_imag[135] = 16'h15E2;
w_real[136] = 16'h8276; w_imag[136] = 16'h18F8;
w_real[137] = 16'h831D; w_imag[137] = 16'h1C0B;
w_real[138] = 16'h83D7; w_imag[138] = 16'h1F19;
w_real[139] = 16'h84A3; w_imag[139] = 16'h2223;
w_real[140] = 16'h8583; w_imag[140] = 16'h2528;
w_real[141] = 16'h8676; w_imag[141] = 16'h2826;
w_real[142] = 16'h877C; w_imag[142] = 16'h2B1F;
w_real[143] = 16'h8894; w_imag[143] = 16'h2E11;
w_real[144] = 16'h89BF; w_imag[144] = 16'h30FB;
w_real[145] = 16'h8AFC; w_imag[145] = 16'h33DE;
w_real[146] = 16'h8C4B; w_imag[146] = 16'h36BA;
w_real[147] = 16'h8DAB; w_imag[147] = 16'h398C;
w_real[148] = 16'h8F1E; w_imag[148] = 16'h3C56;
w_real[149] = 16'h90A1; w_imag[149] = 16'h3F17;
w_real[150] = 16'h9236; w_imag[150] = 16'h41CE;
w_real[151] = 16'h93DC; w_imag[151] = 16'h447A;
w_real[152] = 16'h9593; w_imag[152] = 16'h471C;
w_real[153] = 16'h975A; w_imag[153] = 16'h49B4;
w_real[154] = 16'h9931; w_imag[154] = 16'h4C3F;
w_real[155] = 16'h9B18; w_imag[155] = 16'h4EBF;
w_real[156] = 16'h9D0E; w_imag[156] = 16'h5133;
w_real[157] = 16'h9F14; w_imag[157] = 16'h539B;
w_real[158] = 16'hA129; w_imag[158] = 16'h55F5;
w_real[159] = 16'hA34C; w_imag[159] = 16'h5842;
w_real[160] = 16'hA57E; w_imag[160] = 16'h5A82;
w_real[161] = 16'hA7BE; w_imag[161] = 16'h5CB4;
w_real[162] = 16'hAA0B; w_imag[162] = 16'h5ED7;
w_real[163] = 16'hAC65; w_imag[163] = 16'h60EC;
w_real[164] = 16'hAECD; w_imag[164] = 16'h62F2;
w_real[165] = 16'hB141; w_imag[165] = 16'h64E8;
w_real[166] = 16'hB3C1; w_imag[166] = 16'h66CF;
w_real[167] = 16'hB64C; w_imag[167] = 16'h68A6;
w_real[168] = 16'hB8E4; w_imag[168] = 16'h6A6D;
w_real[169] = 16'hBB86; w_imag[169] = 16'h6C24;
w_real[170] = 16'hBE32; w_imag[170] = 16'h6DCA;
w_real[171] = 16'hC0E9; w_imag[171] = 16'h6F5F;
w_real[172] = 16'hC3AA; w_imag[172] = 16'h70E2;
w_real[173] = 16'hC674; w_imag[173] = 16'h7255;
w_real[174] = 16'hC946; w_imag[174] = 16'h73B5;
w_real[175] = 16'hCC22; w_imag[175] = 16'h7504;
w_real[176] = 16'hCF05; w_imag[176] = 16'h7641;
w_real[177] = 16'hD1EF; w_imag[177] = 16'h776C;
w_real[178] = 16'hD4E1; w_imag[178] = 16'h7884;
w_real[179] = 16'hD7DA; w_imag[179] = 16'h798A;
w_real[180] = 16'hDAD8; w_imag[180] = 16'h7A7D;
w_real[181] = 16'hDDDD; w_imag[181] = 16'h7B5D;
w_real[182] = 16'hE0E7; w_imag[182] = 16'h7C29;
w_real[183] = 16'hE3F5; w_imag[183] = 16'h7CE3;
w_real[184] = 16'hE708; w_imag[184] = 16'h7D8A;
w_real[185] = 16'hEA1E; w_imag[185] = 16'h7E1D;
w_real[186] = 16'hED38; w_imag[186] = 16'h7E9D;
w_real[187] = 16'hF055; w_imag[187] = 16'h7F09;
w_real[188] = 16'hF375; w_imag[188] = 16'h7F62;
w_real[189] = 16'hF696; w_imag[189] = 16'h7FA7;
w_real[190] = 16'hF9B9; w_imag[190] = 16'h7FD8;
w_real[191] = 16'hFCDC; w_imag[191] = 16'h7FF6;
w_real[192] = 16'h0000; w_imag[192] = 16'h7FFF;
w_real[193] = 16'h0324; w_imag[193] = 16'h7FF6;
w_real[194] = 16'h0647; w_imag[194] = 16'h7FD8;
w_real[195] = 16'h096A; w_imag[195] = 16'h7FA7;
w_real[196] = 16'h0C8B; w_imag[196] = 16'h7F62;
w_real[197] = 16'h0FAB; w_imag[197] = 16'h7F09;
w_real[198] = 16'h12C8; w_imag[198] = 16'h7E9D;
w_real[199] = 16'h15E2; w_imag[199] = 16'h7E1D;
w_real[200] = 16'h18F8; w_imag[200] = 16'h7D8A;
w_real[201] = 16'h1C0B; w_imag[201] = 16'h7CE3;
w_real[202] = 16'h1F19; w_imag[202] = 16'h7C29;
w_real[203] = 16'h2223; w_imag[203] = 16'h7B5D;
w_real[204] = 16'h2528; w_imag[204] = 16'h7A7D;
w_real[205] = 16'h2826; w_imag[205] = 16'h798A;
w_real[206] = 16'h2B1F; w_imag[206] = 16'h7884;
w_real[207] = 16'h2E11; w_imag[207] = 16'h776C;
w_real[208] = 16'h30FB; w_imag[208] = 16'h7641;
w_real[209] = 16'h33DE; w_imag[209] = 16'h7504;
w_real[210] = 16'h36BA; w_imag[210] = 16'h73B5;
w_real[211] = 16'h398C; w_imag[211] = 16'h7255;
w_real[212] = 16'h3C56; w_imag[212] = 16'h70E2;
w_real[213] = 16'h3F17; w_imag[213] = 16'h6F5F;
w_real[214] = 16'h41CE; w_imag[214] = 16'h6DCA;
w_real[215] = 16'h447A; w_imag[215] = 16'h6C24;
w_real[216] = 16'h471C; w_imag[216] = 16'h6A6D;
w_real[217] = 16'h49B4; w_imag[217] = 16'h68A6;
w_real[218] = 16'h4C3F; w_imag[218] = 16'h66CF;
w_real[219] = 16'h4EBF; w_imag[219] = 16'h64E8;
w_real[220] = 16'h5133; w_imag[220] = 16'h62F2;
w_real[221] = 16'h539B; w_imag[221] = 16'h60EC;
w_real[222] = 16'h55F5; w_imag[222] = 16'h5ED7;
w_real[223] = 16'h5842; w_imag[223] = 16'h5CB4;
w_real[224] = 16'h5A82; w_imag[224] = 16'h5A82;
w_real[225] = 16'h5CB4; w_imag[225] = 16'h5842;
w_real[226] = 16'h5ED7; w_imag[226] = 16'h55F5;
w_real[227] = 16'h60EC; w_imag[227] = 16'h539B;
w_real[228] = 16'h62F2; w_imag[228] = 16'h5133;
w_real[229] = 16'h64E8; w_imag[229] = 16'h4EBF;
w_real[230] = 16'h66CF; w_imag[230] = 16'h4C3F;
w_real[231] = 16'h68A6; w_imag[231] = 16'h49B4;
w_real[232] = 16'h6A6D; w_imag[232] = 16'h471C;
w_real[233] = 16'h6C24; w_imag[233] = 16'h447A;
w_real[234] = 16'h6DCA; w_imag[234] = 16'h41CE;
w_real[235] = 16'h6F5F; w_imag[235] = 16'h3F17;
w_real[236] = 16'h70E2; w_imag[236] = 16'h3C56;
w_real[237] = 16'h7255; w_imag[237] = 16'h398C;
w_real[238] = 16'h73B5; w_imag[238] = 16'h36BA;
w_real[239] = 16'h7504; w_imag[239] = 16'h33DE;
w_real[240] = 16'h7641; w_imag[240] = 16'h30FB;
w_real[241] = 16'h776C; w_imag[241] = 16'h2E11;
w_real[242] = 16'h7884; w_imag[242] = 16'h2B1F;
w_real[243] = 16'h798A; w_imag[243] = 16'h2826;
w_real[244] = 16'h7A7D; w_imag[244] = 16'h2528;
w_real[245] = 16'h7B5D; w_imag[245] = 16'h2223;
w_real[246] = 16'h7C29; w_imag[246] = 16'h1F19;
w_real[247] = 16'h7CE3; w_imag[247] = 16'h1C0B;
w_real[248] = 16'h7D8A; w_imag[248] = 16'h18F8;
w_real[249] = 16'h7E1D; w_imag[249] = 16'h15E2;
w_real[250] = 16'h7E9D; w_imag[250] = 16'h12C8;
w_real[251] = 16'h7F09; w_imag[251] = 16'h0FAB;
w_real[252] = 16'h7F62; w_imag[252] = 16'h0C8B;
w_real[253] = 16'h7FA7; w_imag[253] = 16'h096A;
w_real[254] = 16'h7FD8; w_imag[254] = 16'h0647;
w_real[255] = 16'h7FF6; w_imag[255] = 16'h0324;
