0 0
5 -28
33 -81
136 -203
424 -424
-170 113
-189 78
-163 32
-152 0
-163 -32
-189 -78
-170 -113
424 424
136 203
33 81
5 28
