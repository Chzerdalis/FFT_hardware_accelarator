w_real[0] = 8'h7F; w_imag[0] = 8'h00;
w_real[1] = 8'h7F; w_imag[1] = 8'hF4;
w_real[2] = 8'h7D; w_imag[2] = 8'hE8;
w_real[3] = 8'h7A; w_imag[3] = 8'hDB;
w_real[4] = 8'h76; w_imag[4] = 8'hD0;
w_real[5] = 8'h70; w_imag[5] = 8'hC4;
w_real[6] = 8'h6A; w_imag[6] = 8'hB9;
w_real[7] = 8'h62; w_imag[7] = 8'hAF;
w_real[8] = 8'h5A; w_imag[8] = 8'hA6;
w_real[9] = 8'h51; w_imag[9] = 8'h9E;
w_real[10] = 8'h47; w_imag[10] = 8'h96;
w_real[11] = 8'h3C; w_imag[11] = 8'h90;
w_real[12] = 8'h30; w_imag[12] = 8'h8A;
w_real[13] = 8'h25; w_imag[13] = 8'h86;
w_real[14] = 8'h18; w_imag[14] = 8'h83;
w_real[15] = 8'h0C; w_imag[15] = 8'h81;
w_real[16] = 8'h00; w_imag[16] = 8'h80;
w_real[17] = 8'hF4; w_imag[17] = 8'h81;
w_real[18] = 8'hE8; w_imag[18] = 8'h83;
w_real[19] = 8'hDB; w_imag[19] = 8'h86;
w_real[20] = 8'hD0; w_imag[20] = 8'h8A;
w_real[21] = 8'hC4; w_imag[21] = 8'h90;
w_real[22] = 8'hB9; w_imag[22] = 8'h96;
w_real[23] = 8'hAF; w_imag[23] = 8'h9E;
w_real[24] = 8'hA6; w_imag[24] = 8'hA6;
w_real[25] = 8'h9E; w_imag[25] = 8'hAF;
w_real[26] = 8'h96; w_imag[26] = 8'hB9;
w_real[27] = 8'h90; w_imag[27] = 8'hC4;
w_real[28] = 8'h8A; w_imag[28] = 8'hD0;
w_real[29] = 8'h86; w_imag[29] = 8'hDB;
w_real[30] = 8'h83; w_imag[30] = 8'hE8;
w_real[31] = 8'h81; w_imag[31] = 8'hF4;
w_real[32] = 8'h80; w_imag[32] = 8'h00;
w_real[33] = 8'h81; w_imag[33] = 8'h0C;
w_real[34] = 8'h83; w_imag[34] = 8'h18;
w_real[35] = 8'h86; w_imag[35] = 8'h25;
w_real[36] = 8'h8A; w_imag[36] = 8'h30;
w_real[37] = 8'h90; w_imag[37] = 8'h3C;
w_real[38] = 8'h96; w_imag[38] = 8'h47;
w_real[39] = 8'h9E; w_imag[39] = 8'h51;
w_real[40] = 8'hA6; w_imag[40] = 8'h5A;
w_real[41] = 8'hAF; w_imag[41] = 8'h62;
w_real[42] = 8'hB9; w_imag[42] = 8'h6A;
w_real[43] = 8'hC4; w_imag[43] = 8'h70;
w_real[44] = 8'hD0; w_imag[44] = 8'h76;
w_real[45] = 8'hDB; w_imag[45] = 8'h7A;
w_real[46] = 8'hE8; w_imag[46] = 8'h7D;
w_real[47] = 8'hF4; w_imag[47] = 8'h7F;
w_real[48] = 8'h00; w_imag[48] = 8'h7F;
w_real[49] = 8'h0C; w_imag[49] = 8'h7F;
w_real[50] = 8'h18; w_imag[50] = 8'h7D;
w_real[51] = 8'h25; w_imag[51] = 8'h7A;
w_real[52] = 8'h30; w_imag[52] = 8'h76;
w_real[53] = 8'h3C; w_imag[53] = 8'h70;
w_real[54] = 8'h47; w_imag[54] = 8'h6A;
w_real[55] = 8'h51; w_imag[55] = 8'h62;
w_real[56] = 8'h5A; w_imag[56] = 8'h5A;
w_real[57] = 8'h62; w_imag[57] = 8'h51;
w_real[58] = 8'h6A; w_imag[58] = 8'h47;
w_real[59] = 8'h70; w_imag[59] = 8'h3C;
w_real[60] = 8'h76; w_imag[60] = 8'h30;
w_real[61] = 8'h7A; w_imag[61] = 8'h25;
w_real[62] = 8'h7D; w_imag[62] = 8'h18;
w_real[63] = 8'h7F; w_imag[63] = 8'h0C;
