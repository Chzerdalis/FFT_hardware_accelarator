gen_input_real[0] = 32'sd0;
gen_input_real[1] = 32'sd32767;
gen_input_real[2] = -32'sd609;
gen_input_real[3] = -32'sd26021;
gen_input_real[4] = 32'sd1595;
gen_input_real[5] = 32'sd19510;
gen_input_real[6] = -32'sd2729;
gen_input_real[7] = -32'sd15929;
gen_input_real[8] = 32'sd3910;
gen_input_real[9] = 32'sd13024;
gen_input_real[10] = -32'sd5655;
gen_input_real[11] = -32'sd9141;
gen_input_real[12] = 32'sd7846;
gen_input_real[13] = 32'sd6167;
gen_input_real[14] = -32'sd9500;
gen_input_real[15] = -32'sd7089;
gen_input_real[16] = 32'sd9488;
gen_input_real[17] = 32'sd10326;
gen_input_real[18] = -32'sd8186;
gen_input_real[19] = -32'sd11345;
gen_input_real[20] = 32'sd7997;
gen_input_real[21] = 32'sd7976;
gen_input_real[22] = -32'sd9273;
gen_input_real[23] = -32'sd1727;
gen_input_real[24] = 32'sd9925;
gen_input_real[25] = -32'sd3975;
gen_input_real[26] = -32'sd9835;
gen_input_real[27] = 32'sd8019;
gen_input_real[28] = 32'sd10199;
gen_input_real[29] = -32'sd11693;
gen_input_real[30] = -32'sd11091;
gen_input_real[31] = 32'sd14416;
gen_input_real[32] = 32'sd11988;
gen_input_real[33] = -32'sd13998;
gen_input_real[34] = -32'sd12181;
gen_input_real[35] = 32'sd9912;
gen_input_real[36] = 32'sd11092;
gen_input_real[37] = -32'sd4816;
gen_input_real[38] = -32'sd9045;
gen_input_real[39] = 32'sd1870;
gen_input_real[40] = 32'sd7881;
gen_input_real[41] = -32'sd960;
gen_input_real[42] = -32'sd8876;
gen_input_real[43] = 32'sd981;
gen_input_real[44] = 32'sd10036;
gen_input_real[45] = -32'sd2148;
gen_input_real[46] = -32'sd9601;
gen_input_real[47] = 32'sd4378;
gen_input_real[48] = 32'sd8752;
gen_input_real[49] = -32'sd6791;
gen_input_real[50] = -32'sd8600;
gen_input_real[51] = 32'sd7467;
gen_input_real[52] = 32'sd8475;
gen_input_real[53] = -32'sd5095;
gen_input_real[54] = -32'sd6795;
gen_input_real[55] = 32'sd1691;
gen_input_real[56] = 32'sd3832;
gen_input_real[57] = 32'sd376;
gen_input_real[58] = -32'sd1674;
gen_input_real[59] = -32'sd2009;
gen_input_real[60] = 32'sd653;
gen_input_real[61] = 32'sd4037;
gen_input_real[62] = -32'sd341;
gen_input_real[63] = -32'sd4453;
gen_input_real[64] = 32'sd875;
gen_input_real[65] = 32'sd1931;
gen_input_real[66] = -32'sd1192;
gen_input_real[67] = 32'sd1810;
gen_input_real[68] = 32'sd589;
gen_input_real[69] = -32'sd4431;
gen_input_real[70] = 32'sd374;
gen_input_real[71] = 32'sd5559;
gen_input_real[72] = -32'sd1745;
gen_input_real[73] = -32'sd5947;
gen_input_real[74] = 32'sd3476;
gen_input_real[75] = 32'sd5442;
gen_input_real[76] = -32'sd4925;
gen_input_real[77] = -32'sd3857;
gen_input_real[78] = 32'sd5750;
gen_input_real[79] = 32'sd2133;
gen_input_real[80] = -32'sd5403;
gen_input_real[81] = -32'sd792;
gen_input_real[82] = 32'sd3434;
gen_input_real[83] = -32'sd351;
gen_input_real[84] = -32'sd532;
gen_input_real[85] = 32'sd500;
gen_input_real[86] = -32'sd2004;
gen_input_real[87] = 32'sd1075;
gen_input_real[88] = 32'sd3657;
gen_input_real[89] = -32'sd3291;
gen_input_real[90] = -32'sd4571;
gen_input_real[91] = 32'sd4840;
gen_input_real[92] = 32'sd4339;
gen_input_real[93] = -32'sd5620;
gen_input_real[94] = -32'sd3003;
gen_input_real[95] = 32'sd5607;
gen_input_real[96] = 32'sd2161;
gen_input_real[97] = -32'sd4811;
gen_input_real[98] = -32'sd2944;
gen_input_real[99] = 32'sd4203;
gen_input_real[100] = 32'sd4408;
gen_input_real[101] = -32'sd3927;
gen_input_real[102] = -32'sd5486;
gen_input_real[103] = 32'sd2978;
gen_input_real[104] = 32'sd6757;
gen_input_real[105] = -32'sd2013;
gen_input_real[106] = -32'sd8781;
gen_input_real[107] = 32'sd2948;
gen_input_real[108] = 32'sd9985;
gen_input_real[109] = -32'sd6257;
gen_input_real[110] = -32'sd8370;
gen_input_real[111] = 32'sd10089;
gen_input_real[112] = 32'sd4647;
gen_input_real[113] = -32'sd12025;
gen_input_real[114] = -32'sd728;
gen_input_real[115] = 32'sd12023;
gen_input_real[116] = -32'sd2476;
gen_input_real[117] = -32'sd12135;
gen_input_real[118] = 32'sd4149;
gen_input_real[119] = 32'sd12914;
gen_input_real[120] = -32'sd4742;
gen_input_real[121] = -32'sd12215;
gen_input_real[122] = 32'sd5909;
gen_input_real[123] = 32'sd8806;
gen_input_real[124] = -32'sd6892;
gen_input_real[125] = -32'sd5075;
gen_input_real[126] = 32'sd5852;
gen_input_real[127] = 32'sd4183;
gen_input_real[128] = -32'sd4183;
gen_input_real[129] = -32'sd5852;
gen_input_real[130] = 32'sd5075;
gen_input_real[131] = 32'sd6892;
gen_input_real[132] = -32'sd8806;
gen_input_real[133] = -32'sd5909;
gen_input_real[134] = 32'sd12215;
gen_input_real[135] = 32'sd4742;
gen_input_real[136] = -32'sd12914;
gen_input_real[137] = -32'sd4149;
gen_input_real[138] = 32'sd12135;
gen_input_real[139] = 32'sd2476;
gen_input_real[140] = -32'sd12023;
gen_input_real[141] = 32'sd728;
gen_input_real[142] = 32'sd12025;
gen_input_real[143] = -32'sd4647;
gen_input_real[144] = -32'sd10089;
gen_input_real[145] = 32'sd8370;
gen_input_real[146] = 32'sd6257;
gen_input_real[147] = -32'sd9985;
gen_input_real[148] = -32'sd2948;
gen_input_real[149] = 32'sd8781;
gen_input_real[150] = 32'sd2013;
gen_input_real[151] = -32'sd6757;
gen_input_real[152] = -32'sd2978;
gen_input_real[153] = 32'sd5486;
gen_input_real[154] = 32'sd3927;
gen_input_real[155] = -32'sd4408;
gen_input_real[156] = -32'sd4203;
gen_input_real[157] = 32'sd2944;
gen_input_real[158] = 32'sd4811;
gen_input_real[159] = -32'sd2161;
gen_input_real[160] = -32'sd5607;
gen_input_real[161] = 32'sd3003;
gen_input_real[162] = 32'sd5620;
gen_input_real[163] = -32'sd4339;
gen_input_real[164] = -32'sd4840;
gen_input_real[165] = 32'sd4571;
gen_input_real[166] = 32'sd3291;
gen_input_real[167] = -32'sd3657;
gen_input_real[168] = -32'sd1075;
gen_input_real[169] = 32'sd2004;
gen_input_real[170] = -32'sd500;
gen_input_real[171] = 32'sd532;
gen_input_real[172] = 32'sd351;
gen_input_real[173] = -32'sd3434;
gen_input_real[174] = 32'sd792;
gen_input_real[175] = 32'sd5403;
gen_input_real[176] = -32'sd2133;
gen_input_real[177] = -32'sd5750;
gen_input_real[178] = 32'sd3857;
gen_input_real[179] = 32'sd4925;
gen_input_real[180] = -32'sd5442;
gen_input_real[181] = -32'sd3476;
gen_input_real[182] = 32'sd5947;
gen_input_real[183] = 32'sd1745;
gen_input_real[184] = -32'sd5559;
gen_input_real[185] = -32'sd374;
gen_input_real[186] = 32'sd4431;
gen_input_real[187] = -32'sd589;
gen_input_real[188] = -32'sd1810;
gen_input_real[189] = 32'sd1192;
gen_input_real[190] = -32'sd1931;
gen_input_real[191] = -32'sd875;
gen_input_real[192] = 32'sd4453;
gen_input_real[193] = 32'sd341;
gen_input_real[194] = -32'sd4037;
gen_input_real[195] = -32'sd653;
gen_input_real[196] = 32'sd2009;
gen_input_real[197] = 32'sd1674;
gen_input_real[198] = -32'sd376;
gen_input_real[199] = -32'sd3832;
gen_input_real[200] = -32'sd1691;
gen_input_real[201] = 32'sd6795;
gen_input_real[202] = 32'sd5095;
gen_input_real[203] = -32'sd8475;
gen_input_real[204] = -32'sd7467;
gen_input_real[205] = 32'sd8600;
gen_input_real[206] = 32'sd6791;
gen_input_real[207] = -32'sd8752;
gen_input_real[208] = -32'sd4378;
gen_input_real[209] = 32'sd9601;
gen_input_real[210] = 32'sd2148;
gen_input_real[211] = -32'sd10036;
gen_input_real[212] = -32'sd981;
gen_input_real[213] = 32'sd8876;
gen_input_real[214] = 32'sd960;
gen_input_real[215] = -32'sd7881;
gen_input_real[216] = -32'sd1870;
gen_input_real[217] = 32'sd9045;
gen_input_real[218] = 32'sd4816;
gen_input_real[219] = -32'sd11092;
gen_input_real[220] = -32'sd9912;
gen_input_real[221] = 32'sd12181;
gen_input_real[222] = 32'sd13998;
gen_input_real[223] = -32'sd11988;
gen_input_real[224] = -32'sd14416;
gen_input_real[225] = 32'sd11091;
gen_input_real[226] = 32'sd11693;
gen_input_real[227] = -32'sd10199;
gen_input_real[228] = -32'sd8019;
gen_input_real[229] = 32'sd9835;
gen_input_real[230] = 32'sd3975;
gen_input_real[231] = -32'sd9925;
gen_input_real[232] = 32'sd1727;
gen_input_real[233] = 32'sd9273;
gen_input_real[234] = -32'sd7976;
gen_input_real[235] = -32'sd7997;
gen_input_real[236] = 32'sd11345;
gen_input_real[237] = 32'sd8186;
gen_input_real[238] = -32'sd10326;
gen_input_real[239] = -32'sd9488;
gen_input_real[240] = 32'sd7089;
gen_input_real[241] = 32'sd9500;
gen_input_real[242] = -32'sd6167;
gen_input_real[243] = -32'sd7846;
gen_input_real[244] = 32'sd9141;
gen_input_real[245] = 32'sd5655;
gen_input_real[246] = -32'sd13024;
gen_input_real[247] = -32'sd3910;
gen_input_real[248] = 32'sd15929;
gen_input_real[249] = 32'sd2729;
gen_input_real[250] = -32'sd19510;
gen_input_real[251] = -32'sd1595;
gen_input_real[252] = 32'sd26021;
gen_input_real[253] = 32'sd609;
gen_input_real[254] = -32'sd32767;
gen_input_real[255] = 32'sd0;
