gen_input_real[0] = 18'sd0;
gen_input_real[16] = 18'sd255;
gen_input_real[32] = 18'sd15;
gen_input_real[48] = -18'sd183;
gen_input_real[4] = -18'sd34;
gen_input_real[20] = 18'sd114;
gen_input_real[36] = 18'sd31;
gen_input_real[52] = -18'sd73;
gen_input_real[8] = 18'sd13;
gen_input_real[24] = 18'sd45;
gen_input_real[40] = -18'sd66;
gen_input_real[56] = -18'sd23;
gen_input_real[12] = 18'sd72;
gen_input_real[28] = 18'sd11;
gen_input_real[44] = -18'sd35;
gen_input_real[60] = -18'sd7;
gen_input_real[1] = 18'sd3;
gen_input_real[17] = -18'sd10;
gen_input_real[33] = 18'sd9;
gen_input_real[49] = 18'sd45;
gen_input_real[5] = -18'sd12;
gen_input_real[21] = -18'sd72;
gen_input_real[37] = 18'sd0;
gen_input_real[53] = 18'sd76;
gen_input_real[9] = 18'sd24;
gen_input_real[25] = -18'sd58;
gen_input_real[41] = -18'sd38;
gen_input_real[57] = 18'sd30;
gen_input_real[13] = 18'sd39;
gen_input_real[29] = -18'sd2;
gen_input_real[45] = -18'sd37;
gen_input_real[61] = -18'sd23;
gen_input_real[2] = 18'sd23;
gen_input_real[18] = 18'sd37;
gen_input_real[34] = 18'sd2;
gen_input_real[50] = -18'sd39;
gen_input_real[6] = -18'sd30;
gen_input_real[22] = 18'sd38;
gen_input_real[38] = 18'sd58;
gen_input_real[54] = -18'sd24;
gen_input_real[10] = -18'sd76;
gen_input_real[26] = 18'sd0;
gen_input_real[42] = 18'sd72;
gen_input_real[58] = 18'sd12;
gen_input_real[14] = -18'sd45;
gen_input_real[30] = -18'sd9;
gen_input_real[46] = 18'sd10;
gen_input_real[62] = -18'sd3;
gen_input_real[3] = 18'sd7;
gen_input_real[19] = 18'sd35;
gen_input_real[35] = -18'sd11;
gen_input_real[51] = -18'sd72;
gen_input_real[7] = 18'sd23;
gen_input_real[23] = 18'sd66;
gen_input_real[39] = -18'sd45;
gen_input_real[55] = -18'sd13;
gen_input_real[11] = 18'sd73;
gen_input_real[27] = -18'sd31;
gen_input_real[43] = -18'sd114;
gen_input_real[59] = 18'sd34;
gen_input_real[15] = 18'sd183;
gen_input_real[31] = -18'sd15;
gen_input_real[47] = -18'sd255;
gen_input_real[63] = 18'sd0;
