0 0
0 -115
1 -217
3 -332
5 -452
8 -548
12 -682
16 -788
22 -900
27 -1011
34 -1127
42 -1256
50 -1360
58 -1461
68 -1588
78 -1703
88 -1807
100 -1922
111 -2019
125 -2152
138 -2256
153 -2375
169 -2500
182 -2587
199 -2709
218 -2848
236 -2961
255 -3077
274 -3190
295 -3315
319 -3460
339 -3562
362 -3680
386 -3806
411 -3930
438 -4064
463 -4177
489 -4296
519 -4432
550 -4576
586 -4754
862 -6817
637 -4919
980 -7387
682 -5025
724 -5211
762 -5366
800 -5512
839 -5660
876 -5786
921 -5960
962 -6098
1003 -6237
1046 -6379
1096 -6555
1142 -6707
1194 -6886
1250 -7078
1312 -7296
1389 -7591
1505 -8087
3341 -17644
3320 -17247
1319 -6742
1464 -7363
1552 -7683
1630 -7941
1703 -8170
1780 -8408
1860 -8658
1952 -8950
2064 -9326
2277 -10143
6517 -28614
1774 -7681
2020 -8625
2145 -9035
2251 -9353
2345 -9612
2430 -9832
2522 -10071
2607 -10277
2689 -10464
2779 -10680
2869 -10888
2969 -11127
3060 -11328
3173 -11604
3262 -11788
3368 -12029
3471 -12253
3587 -12515
3707 -12785
3830 -13057
3958 -13344
4088 -13628
4228 -13939
4383 -14291
4547 -14666
4716 -15048
4912 -15505
5119 -15989
5368 -16591
5656 -17299
6013 -18203
6506 -19494
7281 -21595
9032 -26518
37605 -109312
3638 -10470
7416 -21134
40301 -113735
941 -2632
3687 -10207
4829 -13240
5683 -15435
6555 -17634
7778 -20730
10534 -27818
55665 -145636
-748 1940
2993 -7689
4313 -10981
5069 -12791
5622 -14058
6073 -15053
6463 -15880
6828 -16628
7167 -17304
7515 -17987
7865 -18665
8214 -19326
8580 -20016
8959 -20726
9375 -21505
9823 -22345
10323 -23289
10904 -24397
11575 -25688
12424 -27347
13538 -29556
15216 -32953
18196 -39091
25839 -55068
137699 -291141
-10032 21045
1532 -3188
5280 -10903
7312 -14982
8674 -17634
9774 -19719
10693 -21408
11558 -22963
12404 -24456
13266 -25957
14155 -27488
15142 -29185
16254 -31095
17594 -33408
19252 -36285
21492 -40209
24878 -46202
30962 -57081
46736 -85535
253242 -460112
-30902 55739
-5568 9972
2351 -4180
6457 -11398
9130 -16003
11148 -19401
12818 -22150
14266 -24479
15636 -26640
16941 -28662
18245 -30653
19595 -32692
21024 -34835
22534 -37077
24233 -39599
26150 -42438
28384 -45750
31143 -49855
34642 -55079
39466 -62324
46793 -73395
59975 -93438
93835 -145208
484048 -744035
-78823 120351
-20268 30739
-2042 3077
7756 -11608
14639 -21764
20387 -30109
25977 -38114
32111 -46803
39760 -57574
50769 -73035
70059 -100127
118853 -168759
649274 -915917
-137052 192085
-49878 69454
-23867 33020
-10815 14867
-2579 3523
3373 -4577
8121 -10950
12122 -16241
15711 -20914
19095 -25258
22368 -29399
25647 -33495
29106 -37771
32759 -42243
36810 -47168
41432 -52756
46908 -59353
53621 -67420
62375 -77935
74569 -92587
93506 -115374
128123 -157099
217083 -264516
1100966 -1333170
-277114 333471
-104867 125410
-55173 65571
-30727 36292
-15562 18266
-4764 5557
3611 -4186
10668 -12291
16906 -19357
22681 -25810
28228 -31924
33769 -37955
39442 -44058
45376 -50375
51745 -57092
58746 -64418
66621 -72604
75675 -81966
86339 -92943
99236 -106171
115393 -122700
136543 -144300
165813 -174158
210063 -219285
287276 -298052
469942 -484585
1965078 -2013910
-381365 388451
129234 -130830
1760247 -1771081
-752487 752487
-361727 359514
-244349 241369
-184752 181382
-147476 143900
-121282 117617
-101453 97785
-85488 81893
-72007 68556
-60117 56886
-49137 46211
-38528 36011
-27787 25813
-16319 15067
-3286 3015
12572 -11465
33685 -30530
65291 -58813
121599 -108860
261880 -233000
1421789 -1257202
-588514 517178
-272451 237949
-186386 161778
-145522 125528
-121088 103805
-104589 89105
-92508 78325
-83130 69947
-75493 63127
-69122 57440
-63596 52519
-58716 48187
-54316 44297
-50248 40724
-46443 37405
-42875 34315
-39351 31296
-35860 28341
-32407 25451
-28816 22488
-25107 19470
-21096 16256
-16725 12806
-11731 8926
-5934 4486
1200 -902
10413 -7772
23209 -17213
42862 -31585
78326 -57349
166196 -120905
828855 -599096
-400897 287900
-181368 129405
-123485 87535
-96181 67738
-79856 55875
-68742 47785
-60436 41737
-53880 36966
-48413 32997
-43641 29549
-39315 26444
-35332 23608
-31498 20906
-27753 18298
-23978 15704
-20045 13041
-15837 10234
-11277 7238
-6083 3878
0 0
7555 -4752
17531 -10951
32076 -19901
56859 -35035
114529 -70087
504036 -306327
-250350 151100
-96520 57851
-51991 30945
-25397 15011
-1785 1047
27758 -16177
84255 -48759
416331 -239235
-211425 120629
-59944 33958
20522 -11542
333567 -186269
-237693 131776
-99432 54726
-44451 24288
18636 -10109
301513 -162353
-180877 96681
178714 -94821
-292026 153795
-171094 89436
-134906 69994
-115698 59578
-103158 52721
-94027 47691
-86848 43715
-80927 40424
-75793 37570
-71142 34993
-66744 32575
-62384 30211
-57732 27740
-52322 24943
-45250 21402
-34071 15987
-9338 4346
142345 -65728
-177050 81094
-104589 47518
-86059 38781
-77030 34428
-71384 31642
-67315 29592
-64131 27958
-61457 26568
-59113 25339
-56980 24219
-54897 23135
-52898 22101
-50833 21055
-48607 19959
-46085 18758
-42985 17343
-38807 15519
-32139 12738
-17731 6965
64282 -25023
-112945 43567
-67414 25767
-52237 19782
-36160 13567
34444 -12803
-115869 42665
-77429 28241
-67274 24304
-62055 22203
-58523 20737
-55778 19572
-53379 18547
-50935 17522
-48155 16401
-44164 14891
-36057 12034
7835 -2588
-91503 29917
-65836 21302
-59335 18997
-56064 17761
-53869 16884
-52174 16177
-50626 15527
-49152 14910
-47385 14215
-44924 13327
-39897 11702
-13407 3888
-75077 21522
-58582 16599
-54563 15280
-52512 14532
-51245 14012
-50339 13598
-49619 13241
-49009 12917
-48492 12622
-48031 12344
-47626 12085
-47252 11836
-46919 11599
-46590 11366
-46302 11146
-46037 10933
-45757 10718
-45512 10513
-45270 10311
-45057 10118
-44857 9928
-44638 9736
-44432 9549
-44248 9367
-44066 9187
-43889 9010
-43718 8835
-43561 8664
-43403 8495
-43255 8328
-43121 8165
-42988 8003
-42837 7839
-42710 7681
-42569 7521
-42469 7369
-42349 7214
-42229 7060
-42124 6910
-42010 6759
-41907 6611
-41785 6460
-41689 6314
-41605 6171
-41528 6030
-41430 5886
-41339 5743
-41246 5601
-41180 5464
-41099 5325
-41053 5191
-40952 5051
-40903 4917
-40819 4780
-40741 4644
-40682 4511
-40622 4378
-40548 4245
-40511 4115
-40444 3983
-40403 3854
-40323 3721
-40275 3592
-40215 3463
-40173 3335
-40098 3205
-39916 3067
-40252 2969
-40098 2834
-40028 2705
-39996 2580
-39946 2454
-39928 2330
-39885 2204
-39863 2080
-39828 1956
-39792 1832
-39779 1709
-39758 1586
-39738 1463
-39712 1340
-39715 1218
-39680 1095
-39667 973
-39671 852
-39645 729
-39651 608
-39629 486
-39644 364
-39625 243
-39632 121
-39630 0
-39632 -121
-39625 -243
-39644 -364
-39629 -486
-39651 -608
-39645 -729
-39671 -852
-39667 -973
-39680 -1095
-39715 -1218
-39712 -1340
-39738 -1463
-39758 -1586
-39779 -1709
-39792 -1832
-39828 -1956
-39863 -2080
-39885 -2204
-39928 -2330
-39946 -2454
-39996 -2580
-40028 -2705
-40098 -2834
-40252 -2969
-39916 -3067
-40098 -3205
-40173 -3335
-40215 -3463
-40275 -3592
-40323 -3721
-40403 -3854
-40444 -3983
-40511 -4115
-40548 -4245
-40622 -4378
-40682 -4511
-40741 -4644
-40819 -4780
-40903 -4917
-40952 -5051
-41053 -5191
-41099 -5325
-41180 -5464
-41246 -5601
-41339 -5743
-41430 -5886
-41528 -6030
-41605 -6171
-41689 -6314
-41785 -6460
-41907 -6611
-42010 -6759
-42124 -6910
-42229 -7060
-42349 -7214
-42469 -7369
-42569 -7521
-42710 -7681
-42837 -7839
-42988 -8003
-43121 -8165
-43255 -8328
-43403 -8495
-43561 -8664
-43718 -8835
-43889 -9010
-44066 -9187
-44248 -9367
-44432 -9549
-44638 -9736
-44857 -9928
-45057 -10118
-45270 -10311
-45512 -10513
-45757 -10718
-46037 -10933
-46302 -11146
-46590 -11366
-46919 -11599
-47252 -11836
-47626 -12085
-48031 -12344
-48492 -12622
-49009 -12917
-49619 -13241
-50339 -13598
-51245 -14012
-52512 -14532
-54563 -15280
-58582 -16599
-75077 -21522
-13407 -3888
-39897 -11702
-44924 -13327
-47385 -14215
-49152 -14910
-50626 -15527
-52174 -16177
-53869 -16884
-56064 -17761
-59335 -18997
-65836 -21302
-91503 -29917
7835 2588
-36057 -12034
-44164 -14891
-48155 -16401
-50935 -17522
-53379 -18547
-55778 -19572
-58523 -20737
-62055 -22203
-67274 -24304
-77429 -28241
-115869 -42665
34444 12803
-36160 -13567
-52237 -19782
-67414 -25767
-112945 -43567
64282 25023
-17731 -6965
-32139 -12738
-38807 -15519
-42985 -17343
-46085 -18758
-48607 -19959
-50833 -21055
-52898 -22101
-54897 -23135
-56980 -24219
-59113 -25339
-61457 -26568
-64131 -27958
-67315 -29592
-71384 -31642
-77030 -34428
-86059 -38781
-104589 -47518
-177050 -81094
142345 65728
-9338 -4346
-34071 -15987
-45250 -21402
-52322 -24943
-57732 -27740
-62384 -30211
-66744 -32575
-71142 -34993
-75793 -37570
-80927 -40424
-86848 -43715
-94027 -47691
-103158 -52721
-115698 -59578
-134906 -69994
-171094 -89436
-292026 -153795
178714 94821
-180877 -96681
301513 162353
18636 10109
-44451 -24288
-99432 -54726
-237693 -131776
333567 186269
20522 11542
-59944 -33958
-211425 -120629
416331 239235
84255 48759
27758 16177
-1785 -1047
-25397 -15011
-51991 -30945
-96520 -57851
-250350 -151100
504036 306327
114529 70087
56859 35035
32076 19901
17531 10951
7555 4752
0 0
-6083 -3878
-11277 -7238
-15837 -10234
-20045 -13041
-23978 -15704
-27753 -18298
-31498 -20906
-35332 -23608
-39315 -26444
-43641 -29549
-48413 -32997
-53880 -36966
-60436 -41737
-68742 -47785
-79856 -55875
-96181 -67738
-123485 -87535
-181368 -129405
-400897 -287900
828855 599096
166196 120905
78326 57349
42862 31585
23209 17213
10413 7772
1200 902
-5934 -4486
-11731 -8926
-16725 -12806
-21096 -16256
-25107 -19470
-28816 -22488
-32407 -25451
-35860 -28341
-39351 -31296
-42875 -34315
-46443 -37405
-50248 -40724
-54316 -44297
-58716 -48187
-63596 -52519
-69122 -57440
-75493 -63127
-83130 -69947
-92508 -78325
-104589 -89105
-121088 -103805
-145522 -125528
-186386 -161778
-272451 -237949
-588514 -517178
1421789 1257202
261880 233000
121599 108860
65291 58813
33685 30530
12572 11465
-3286 -3015
-16319 -15067
-27787 -25813
-38528 -36011
-49137 -46211
-60117 -56886
-72007 -68556
-85488 -81893
-101453 -97785
-121282 -117617
-147476 -143900
-184752 -181382
-244349 -241369
-361727 -359514
-752487 -752487
1760247 1771081
129234 130830
-381365 -388451
1965078 2013910
469942 484585
287276 298052
210063 219285
165813 174158
136543 144300
115393 122700
99236 106171
86339 92943
75675 81966
66621 72604
58746 64418
51745 57092
45376 50375
39442 44058
33769 37955
28228 31924
22681 25810
16906 19357
10668 12291
3611 4186
-4764 -5557
-15562 -18266
-30727 -36292
-55173 -65571
-104867 -125410
-277114 -333471
1100966 1333170
217083 264516
128123 157099
93506 115374
74569 92587
62375 77935
53621 67420
46908 59353
41432 52756
36810 47168
32759 42243
29106 37771
25647 33495
22368 29399
19095 25258
15711 20914
12122 16241
8121 10950
3373 4577
-2579 -3523
-10815 -14867
-23867 -33020
-49878 -69454
-137052 -192085
649274 915917
118853 168759
70059 100127
50769 73035
39760 57574
32111 46803
25977 38114
20387 30109
14639 21764
7756 11608
-2042 -3077
-20268 -30739
-78823 -120351
484048 744035
93835 145208
59975 93438
46793 73395
39466 62324
34642 55079
31143 49855
28384 45750
26150 42438
24233 39599
22534 37077
21024 34835
19595 32692
18245 30653
16941 28662
15636 26640
14266 24479
12818 22150
11148 19401
9130 16003
6457 11398
2351 4180
-5568 -9972
-30902 -55739
253242 460112
46736 85535
30962 57081
24878 46202
21492 40209
19252 36285
17594 33408
16254 31095
15142 29185
14155 27488
13266 25957
12404 24456
11558 22963
10693 21408
9774 19719
8674 17634
7312 14982
5280 10903
1532 3188
-10032 -21045
137699 291141
25839 55068
18196 39091
15216 32953
13538 29556
12424 27347
11575 25688
10904 24397
10323 23289
9823 22345
9375 21505
8959 20726
8580 20016
8214 19326
7865 18665
7515 17987
7167 17304
6828 16628
6463 15880
6073 15053
5622 14058
5069 12791
4313 10981
2993 7689
-748 -1940
55665 145636
10534 27818
7778 20730
6555 17634
5683 15435
4829 13240
3687 10207
941 2632
40301 113735
7416 21134
3638 10470
37605 109312
9032 26518
7281 21595
6506 19494
6013 18203
5656 17299
5368 16591
5119 15989
4912 15505
4716 15048
4547 14666
4383 14291
4228 13939
4088 13628
3958 13344
3830 13057
3707 12785
3587 12515
3471 12253
3368 12029
3262 11788
3173 11604
3060 11328
2969 11127
2869 10888
2779 10680
2689 10464
2607 10277
2522 10071
2430 9832
2345 9612
2251 9353
2145 9035
2020 8625
1774 7681
6517 28614
2277 10143
2064 9326
1952 8950
1860 8658
1780 8408
1703 8170
1630 7941
1552 7683
1464 7363
1319 6742
3320 17247
3341 17644
1505 8087
1389 7591
1312 7296
1250 7078
1194 6886
1142 6707
1096 6555
1046 6379
1003 6237
962 6098
921 5960
876 5786
839 5660
800 5512
762 5366
724 5211
682 5025
980 7387
637 4919
862 6817
586 4754
550 4576
519 4432
489 4296
463 4177
438 4064
411 3930
386 3806
362 3680
339 3562
319 3460
295 3315
274 3190
255 3077
236 2961
218 2848
199 2709
182 2587
169 2500
153 2375
138 2256
125 2152
111 2019
100 1922
88 1807
78 1703
68 1588
58 1461
50 1360
42 1256
34 1127
27 1011
22 900
16 788
12 682
8 548
5 452
3 332
1 217
0 115
