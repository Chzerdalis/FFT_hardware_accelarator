gen_input_real[0] = 32'sd0;
gen_input_real[256] = 32'sd32767;
gen_input_real[512] = -32'sd2085;
gen_input_real[768] = -32'sd19335;
gen_input_real[64] = 32'sd963;
gen_input_real[320] = 32'sd8653;
gen_input_real[576] = 32'sd2547;
gen_input_real[832] = -32'sd7035;
gen_input_real[128] = -32'sd4174;
gen_input_real[384] = 32'sd9073;
gen_input_real[640] = 32'sd2057;
gen_input_real[896] = -32'sd10725;
gen_input_real[192] = 32'sd2032;
gen_input_real[448] = 32'sd10567;
gen_input_real[704] = -32'sd4364;
gen_input_real[960] = -32'sd7812;
gen_input_real[16] = 32'sd2436;
gen_input_real[272] = 32'sd5221;
gen_input_real[528] = 32'sd1236;
gen_input_real[784] = -32'sd6746;
gen_input_real[80] = -32'sd2951;
gen_input_real[336] = 32'sd9639;
gen_input_real[592] = 32'sd1536;
gen_input_real[848] = -32'sd8359;
gen_input_real[144] = 32'sd2125;
gen_input_real[400] = 32'sd4429;
gen_input_real[656] = -32'sd4015;
gen_input_real[912] = -32'sd2677;
gen_input_real[208] = 32'sd841;
gen_input_real[464] = 32'sd3916;
gen_input_real[720] = 32'sd4629;
gen_input_real[976] = -32'sd7215;
gen_input_real[32] = -32'sd8610;
gen_input_real[288] = 32'sd11915;
gen_input_real[544] = 32'sd11291;
gen_input_real[800] = -32'sd15447;
gen_input_real[96] = -32'sd13278;
gen_input_real[352] = 32'sd14897;
gen_input_real[608] = 32'sd13828;
gen_input_real[864] = -32'sd12014;
gen_input_real[160] = -32'sd12980;
gen_input_real[416] = 32'sd11736;
gen_input_real[672] = 32'sd11578;
gen_input_real[928] = -32'sd13410;
gen_input_real[224] = -32'sd9909;
gen_input_real[480] = 32'sd11486;
gen_input_real[736] = 32'sd9027;
gen_input_real[992] = -32'sd5676;
gen_input_real[48] = -32'sd9771;
gen_input_real[304] = 32'sd1896;
gen_input_real[560] = 32'sd9279;
gen_input_real[816] = -32'sd4224;
gen_input_real[112] = -32'sd5124;
gen_input_real[368] = 32'sd9956;
gen_input_real[624] = 32'sd355;
gen_input_real[880] = -32'sd13556;
gen_input_real[176] = 32'sd552;
gen_input_real[432] = 32'sd13369;
gen_input_real[688] = 32'sd1544;
gen_input_real[944] = -32'sd12016;
gen_input_real[240] = -32'sd2298;
gen_input_real[496] = 32'sd11372;
gen_input_real[752] = 32'sd1478;
gen_input_real[1008] = -32'sd9697;
gen_input_real[4] = -32'sd1261;
gen_input_real[260] = 32'sd6293;
gen_input_real[516] = 32'sd1521;
gen_input_real[772] = -32'sd3003;
gen_input_real[68] = -32'sd2373;
gen_input_real[324] = 32'sd696;
gen_input_real[580] = 32'sd4581;
gen_input_real[836] = -32'sd863;
gen_input_real[132] = -32'sd7539;
gen_input_real[388] = 32'sd3798;
gen_input_real[644] = 32'sd10494;
gen_input_real[900] = -32'sd5640;
gen_input_real[196] = -32'sd13848;
gen_input_real[452] = 32'sd4207;
gen_input_real[708] = 32'sd16469;
gen_input_real[964] = -32'sd1237;
gen_input_real[20] = -32'sd15024;
gen_input_real[276] = -32'sd2287;
gen_input_real[532] = 32'sd10472;
gen_input_real[788] = 32'sd6270;
gen_input_real[84] = -32'sd7124;
gen_input_real[340] = -32'sd8371;
gen_input_real[596] = 32'sd4955;
gen_input_real[852] = 32'sd5422;
gen_input_real[148] = -32'sd4135;
gen_input_real[404] = 32'sd1392;
gen_input_real[660] = 32'sd7784;
gen_input_real[916] = -32'sd7160;
gen_input_real[212] = -32'sd12626;
gen_input_real[468] = 32'sd9790;
gen_input_real[724] = 32'sd12457;
gen_input_real[980] = -32'sd10300;
gen_input_real[36] = -32'sd8743;
gen_input_real[292] = 32'sd9584;
gen_input_real[548] = 32'sd6405;
gen_input_real[804] = -32'sd8256;
gen_input_real[100] = -32'sd6765;
gen_input_real[356] = 32'sd6876;
gen_input_real[612] = 32'sd7734;
gen_input_real[868] = -32'sd6885;
gen_input_real[164] = -32'sd6889;
gen_input_real[420] = 32'sd7577;
gen_input_real[676] = 32'sd3608;
gen_input_real[932] = -32'sd5202;
gen_input_real[228] = -32'sd856;
gen_input_real[484] = 32'sd550;
gen_input_real[740] = 32'sd3719;
gen_input_real[996] = 32'sd2278;
gen_input_real[52] = -32'sd10150;
gen_input_real[308] = -32'sd2637;
gen_input_real[564] = 32'sd11210;
gen_input_real[820] = 32'sd1788;
gen_input_real[116] = -32'sd4739;
gen_input_real[372] = -32'sd1112;
gen_input_real[628] = -32'sd2290;
gen_input_real[884] = 32'sd2464;
gen_input_real[180] = 32'sd4373;
gen_input_real[436] = -32'sd6068;
gen_input_real[692] = -32'sd2814;
gen_input_real[948] = 32'sd9012;
gen_input_real[244] = 32'sd858;
gen_input_real[500] = -32'sd8652;
gen_input_real[756] = 32'sd1033;
gen_input_real[1012] = 32'sd5986;
gen_input_real[8] = -32'sd2792;
gen_input_real[264] = -32'sd3027;
gen_input_real[520] = 32'sd3763;
gen_input_real[776] = -32'sd73;
gen_input_real[72] = -32'sd5455;
gen_input_real[328] = 32'sd3195;
gen_input_real[584] = 32'sd9327;
gen_input_real[840] = -32'sd4542;
gen_input_real[136] = -32'sd13175;
gen_input_real[392] = 32'sd2799;
gen_input_real[648] = 32'sd14036;
gen_input_real[904] = 32'sd441;
gen_input_real[200] = -32'sd11649;
gen_input_real[456] = -32'sd2428;
gen_input_real[712] = 32'sd7464;
gen_input_real[968] = 32'sd2524;
gen_input_real[24] = -32'sd3726;
gen_input_real[280] = -32'sd1567;
gen_input_real[536] = 32'sd2686;
gen_input_real[792] = 32'sd365;
gen_input_real[88] = -32'sd3880;
gen_input_real[344] = 32'sd280;
gen_input_real[600] = 32'sd4643;
gen_input_real[856] = -32'sd717;
gen_input_real[152] = -32'sd4152;
gen_input_real[408] = 32'sd1987;
gen_input_real[664] = 32'sd3143;
gen_input_real[920] = -32'sd3836;
gen_input_real[216] = -32'sd1286;
gen_input_real[472] = 32'sd4464;
gen_input_real[728] = -32'sd3450;
gen_input_real[984] = -32'sd2460;
gen_input_real[40] = 32'sd11455;
gen_input_real[296] = -32'sd669;
gen_input_real[552] = -32'sd16020;
gen_input_real[808] = 32'sd1569;
gen_input_real[104] = 32'sd10997;
gen_input_real[360] = 32'sd1651;
gen_input_real[616] = -32'sd1893;
gen_input_real[872] = -32'sd5951;
gen_input_real[168] = -32'sd2751;
gen_input_real[424] = 32'sd5298;
gen_input_real[680] = 32'sd3136;
gen_input_real[936] = -32'sd28;
gen_input_real[232] = -32'sd3536;
gen_input_real[488] = -32'sd4644;
gen_input_real[744] = 32'sd4006;
gen_input_real[1000] = 32'sd7072;
gen_input_real[56] = -32'sd3099;
gen_input_real[312] = -32'sd6701;
gen_input_real[568] = 32'sd2012;
gen_input_real[824] = 32'sd3668;
gen_input_real[120] = -32'sd496;
gen_input_real[376] = -32'sd2152;
gen_input_real[632] = -32'sd1961;
gen_input_real[888] = 32'sd4436;
gen_input_real[184] = 32'sd1881;
gen_input_real[440] = -32'sd6785;
gen_input_real[696] = 32'sd1420;
gen_input_real[952] = 32'sd5372;
gen_input_real[248] = -32'sd3851;
gen_input_real[504] = -32'sd1032;
gen_input_real[760] = 32'sd4242;
gen_input_real[1016] = -32'sd3505;
gen_input_real[12] = -32'sd3762;
gen_input_real[268] = 32'sd7133;
gen_input_real[524] = 32'sd1911;
gen_input_real[780] = -32'sd9058;
gen_input_real[76] = 32'sd1438;
gen_input_real[332] = 32'sd9289;
gen_input_real[588] = -32'sd3785;
gen_input_real[844] = -32'sd10120;
gen_input_real[140] = 32'sd2515;
gen_input_real[396] = 32'sd11599;
gen_input_real[652] = -32'sd52;
gen_input_real[908] = -32'sd10763;
gen_input_real[204] = 32'sd581;
gen_input_real[460] = 32'sd7159;
gen_input_real[716] = -32'sd1951;
gen_input_real[972] = -32'sd4325;
gen_input_real[28] = -32'sd147;
gen_input_real[284] = 32'sd5575;
gen_input_real[540] = 32'sd3840;
gen_input_real[796] = -32'sd8270;
gen_input_real[92] = -32'sd3888;
gen_input_real[348] = 32'sd6513;
gen_input_real[604] = -32'sd599;
gen_input_real[860] = -32'sd616;
gen_input_real[156] = 32'sd5975;
gen_input_real[412] = -32'sd3625;
gen_input_real[668] = -32'sd9484;
gen_input_real[924] = 32'sd3339;
gen_input_real[220] = 32'sd10564;
gen_input_real[476] = -32'sd250;
gen_input_real[732] = -32'sd9462;
gen_input_real[988] = -32'sd3137;
gen_input_real[44] = 32'sd6916;
gen_input_real[300] = 32'sd5029;
gen_input_real[556] = -32'sd3460;
gen_input_real[812] = -32'sd4254;
gen_input_real[108] = -32'sd705;
gen_input_real[364] = 32'sd2009;
gen_input_real[620] = 32'sd5087;
gen_input_real[876] = -32'sd1559;
gen_input_real[172] = -32'sd8111;
gen_input_real[428] = 32'sd4419;
gen_input_real[684] = 32'sd7670;
gen_input_real[940] = -32'sd8386;
gen_input_real[236] = -32'sd4273;
gen_input_real[492] = 32'sd10566;
gen_input_real[748] = 32'sd1376;
gen_input_real[1004] = -32'sd10516;
gen_input_real[60] = -32'sd1513;
gen_input_real[316] = 32'sd8309;
gen_input_real[572] = 32'sd4813;
gen_input_real[828] = -32'sd5033;
gen_input_real[124] = -32'sd10570;
gen_input_real[380] = 32'sd5084;
gen_input_real[636] = 32'sd15888;
gen_input_real[892] = -32'sd8588;
gen_input_real[188] = -32'sd14576;
gen_input_real[444] = 32'sd8783;
gen_input_real[700] = 32'sd5404;
gen_input_real[956] = -32'sd5132;
gen_input_real[252] = 32'sd3342;
gen_input_real[508] = 32'sd5154;
gen_input_real[764] = -32'sd5401;
gen_input_real[1020] = -32'sd10345;
gen_input_real[1] = 32'sd3307;
gen_input_real[257] = 32'sd14521;
gen_input_real[513] = -32'sd1638;
gen_input_real[769] = -32'sd15184;
gen_input_real[65] = 32'sd2393;
gen_input_real[321] = 32'sd14342;
gen_input_real[577] = -32'sd4169;
gen_input_real[833] = -32'sd11391;
gen_input_real[129] = 32'sd3789;
gen_input_real[385] = 32'sd6816;
gen_input_real[641] = 32'sd24;
gen_input_real[897] = -32'sd5057;
gen_input_real[193] = -32'sd6063;
gen_input_real[449] = 32'sd6400;
gen_input_real[705] = 32'sd10377;
gen_input_real[961] = -32'sd7780;
gen_input_real[17] = -32'sd9104;
gen_input_real[273] = 32'sd8701;
gen_input_real[529] = 32'sd4560;
gen_input_real[785] = -32'sd7551;
gen_input_real[81] = -32'sd2648;
gen_input_real[337] = 32'sd2614;
gen_input_real[593] = 32'sd4970;
gen_input_real[849] = 32'sd2372;
gen_input_real[145] = -32'sd8346;
gen_input_real[401] = -32'sd2647;
gen_input_real[657] = 32'sd10478;
gen_input_real[913] = -32'sd541;
gen_input_real[209] = -32'sd11506;
gen_input_real[465] = 32'sd2052;
gen_input_real[721] = 32'sd10997;
gen_input_real[977] = -32'sd1298;
gen_input_real[33] = -32'sd9964;
gen_input_real[289] = 32'sd2447;
gen_input_real[545] = 32'sd11130;
gen_input_real[801] = -32'sd6056;
gen_input_real[97] = -32'sd12171;
gen_input_real[353] = 32'sd9183;
gen_input_real[609] = 32'sd9103;
gen_input_real[865] = -32'sd11315;
gen_input_real[161] = -32'sd4796;
gen_input_real[417] = 32'sd13625;
gen_input_real[673] = 32'sd4349;
gen_input_real[929] = -32'sd15841;
gen_input_real[225] = -32'sd7917;
gen_input_real[481] = 32'sd16277;
gen_input_real[737] = 32'sd12692;
gen_input_real[993] = -32'sd13351;
gen_input_real[49] = -32'sd16411;
gen_input_real[305] = 32'sd7631;
gen_input_real[561] = 32'sd17185;
gen_input_real[817] = -32'sd3026;
gen_input_real[113] = -32'sd14123;
gen_input_real[369] = 32'sd3031;
gen_input_real[625] = 32'sd9381;
gen_input_real[881] = -32'sd5502;
gen_input_real[177] = -32'sd6284;
gen_input_real[433] = 32'sd6110;
gen_input_real[689] = 32'sd4922;
gen_input_real[945] = -32'sd4823;
gen_input_real[241] = -32'sd3393;
gen_input_real[497] = 32'sd3450;
gen_input_real[753] = 32'sd2481;
gen_input_real[1009] = -32'sd1168;
gen_input_real[5] = -32'sd4090;
gen_input_real[261] = -32'sd2703;
gen_input_real[517] = 32'sd7263;
gen_input_real[773] = 32'sd6111;
gen_input_real[69] = -32'sd9833;
gen_input_real[325] = -32'sd6724;
gen_input_real[581] = 32'sd10388;
gen_input_real[837] = 32'sd3926;
gen_input_real[133] = -32'sd8507;
gen_input_real[389] = 32'sd663;
gen_input_real[645] = 32'sd7084;
gen_input_real[901] = -32'sd4027;
gen_input_real[197] = -32'sd9533;
gen_input_real[453] = 32'sd5177;
gen_input_real[709] = 32'sd13938;
gen_input_real[965] = -32'sd5189;
gen_input_real[21] = -32'sd17243;
gen_input_real[277] = 32'sd3406;
gen_input_real[533] = 32'sd19885;
gen_input_real[789] = 32'sd413;
gen_input_real[85] = -32'sd21128;
gen_input_real[341] = -32'sd3545;
gen_input_real[597] = 32'sd19013;
gen_input_real[853] = 32'sd4268;
gen_input_real[149] = -32'sd16197;
gen_input_real[405] = -32'sd3158;
gen_input_real[661] = 32'sd16626;
gen_input_real[917] = 32'sd1907;
gen_input_real[213] = -32'sd17782;
gen_input_real[469] = -32'sd1590;
gen_input_real[725] = 32'sd15824;
gen_input_real[981] = 32'sd180;
gen_input_real[37] = -32'sd12156;
gen_input_real[293] = 32'sd3518;
gen_input_real[549] = 32'sd7144;
gen_input_real[805] = -32'sd6057;
gen_input_real[101] = -32'sd1106;
gen_input_real[357] = 32'sd3979;
gen_input_real[613] = 32'sd68;
gen_input_real[869] = 32'sd1131;
gen_input_real[165] = -32'sd5576;
gen_input_real[421] = -32'sd4164;
gen_input_real[677] = 32'sd9741;
gen_input_real[933] = 32'sd2563;
gen_input_real[229] = -32'sd8654;
gen_input_real[485] = 32'sd750;
gen_input_real[741] = 32'sd7117;
gen_input_real[997] = -32'sd1076;
gen_input_real[53] = -32'sd7792;
gen_input_real[309] = -32'sd2492;
gen_input_real[565] = 32'sd7787;
gen_input_real[821] = 32'sd5795;
gen_input_real[117] = -32'sd6940;
gen_input_real[373] = -32'sd5754;
gen_input_real[629] = 32'sd8816;
gen_input_real[885] = 32'sd5051;
gen_input_real[181] = -32'sd12151;
gen_input_real[437] = -32'sd6690;
gen_input_real[693] = 32'sd12634;
gen_input_real[949] = 32'sd10409;
gen_input_real[245] = -32'sd11722;
gen_input_real[501] = -32'sd15919;
gen_input_real[757] = 32'sd12351;
gen_input_real[1013] = 32'sd20760;
gen_input_real[9] = -32'sd12465;
gen_input_real[265] = -32'sd19850;
gen_input_real[521] = 32'sd10307;
gen_input_real[777] = 32'sd12818;
gen_input_real[73] = -32'sd8082;
gen_input_real[329] = -32'sd4589;
gen_input_real[585] = 32'sd7378;
gen_input_real[841] = -32'sd779;
gen_input_real[137] = -32'sd7445;
gen_input_real[393] = 32'sd2300;
gen_input_real[649] = 32'sd8644;
gen_input_real[905] = -32'sd348;
gen_input_real[201] = -32'sd10763;
gen_input_real[457] = -32'sd3316;
gen_input_real[713] = 32'sd10664;
gen_input_real[969] = 32'sd5475;
gen_input_real[25] = -32'sd8295;
gen_input_real[281] = -32'sd5086;
gen_input_real[537] = 32'sd8096;
gen_input_real[793] = 32'sd4196;
gen_input_real[89] = -32'sd10514;
gen_input_real[345] = -32'sd3112;
gen_input_real[601] = 32'sd10321;
gen_input_real[857] = 32'sd154;
gen_input_real[153] = -32'sd5892;
gen_input_real[409] = 32'sd1760;
gen_input_real[665] = 32'sd2516;
gen_input_real[921] = 32'sd2061;
gen_input_real[217] = -32'sd4134;
gen_input_real[473] = -32'sd8442;
gen_input_real[729] = 32'sd6881;
gen_input_real[985] = 32'sd11519;
gen_input_real[41] = -32'sd4009;
gen_input_real[297] = -32'sd12329;
gen_input_real[553] = -32'sd3452;
gen_input_real[809] = 32'sd13683;
gen_input_real[105] = 32'sd8031;
gen_input_real[361] = -32'sd14398;
gen_input_real[617] = -32'sd6847;
gen_input_real[873] = 32'sd13843;
gen_input_real[169] = 32'sd2197;
gen_input_real[425] = -32'sd12889;
gen_input_real[681] = 32'sd3127;
gen_input_real[937] = 32'sd9640;
gen_input_real[233] = -32'sd5306;
gen_input_real[489] = -32'sd4054;
gen_input_real[745] = 32'sd2598;
gen_input_real[1001] = 32'sd1857;
gen_input_real[57] = 32'sd426;
gen_input_real[313] = -32'sd5215;
gen_input_real[569] = 32'sd1121;
gen_input_real[825] = 32'sd8996;
gen_input_real[121] = -32'sd6215;
gen_input_real[377] = -32'sd10288;
gen_input_real[633] = 32'sd10842;
gen_input_real[889] = 32'sd10422;
gen_input_real[185] = -32'sd12207;
gen_input_real[441] = -32'sd9660;
gen_input_real[697] = 32'sd9930;
gen_input_real[953] = 32'sd8817;
gen_input_real[249] = -32'sd6042;
gen_input_real[505] = -32'sd8711;
gen_input_real[761] = 32'sd4306;
gen_input_real[1017] = 32'sd7173;
gen_input_real[13] = -32'sd5970;
gen_input_real[269] = -32'sd3262;
gen_input_real[525] = 32'sd6368;
gen_input_real[781] = -32'sd265;
gen_input_real[77] = -32'sd1411;
gen_input_real[333] = 32'sd227;
gen_input_real[589] = -32'sd5354;
gen_input_real[845] = 32'sd3176;
gen_input_real[141] = 32'sd6929;
gen_input_real[397] = -32'sd6371;
gen_input_real[653] = -32'sd3311;
gen_input_real[909] = 32'sd6603;
gen_input_real[205] = 32'sd2587;
gen_input_real[461] = -32'sd4066;
gen_input_real[717] = -32'sd7591;
gen_input_real[973] = 32'sd660;
gen_input_real[29] = 32'sd10877;
gen_input_real[285] = 32'sd1795;
gen_input_real[541] = -32'sd7226;
gen_input_real[797] = -32'sd2811;
gen_input_real[93] = 32'sd241;
gen_input_real[349] = 32'sd2587;
gen_input_real[605] = 32'sd4434;
gen_input_real[861] = -32'sd302;
gen_input_real[157] = -32'sd3845;
gen_input_real[413] = -32'sd4727;
gen_input_real[669] = -32'sd1277;
gen_input_real[925] = 32'sd10861;
gen_input_real[221] = 32'sd5778;
gen_input_real[477] = -32'sd15504;
gen_input_real[733] = -32'sd5078;
gen_input_real[989] = 32'sd16704;
gen_input_real[45] = 32'sd429;
gen_input_real[301] = -32'sd13595;
gen_input_real[557] = 32'sd3103;
gen_input_real[813] = 32'sd7510;
gen_input_real[109] = -32'sd3002;
gen_input_real[365] = -32'sd2514;
gen_input_real[621] = 32'sd1588;
gen_input_real[877] = 32'sd2277;
gen_input_real[173] = -32'sd719;
gen_input_real[429] = -32'sd4880;
gen_input_real[685] = 32'sd149;
gen_input_real[941] = 32'sd5434;
gen_input_real[237] = -32'sd681;
gen_input_real[493] = -32'sd2681;
gen_input_real[749] = 32'sd1732;
gen_input_real[1005] = -32'sd1394;
gen_input_real[61] = 32'sd70;
gen_input_real[317] = 32'sd4282;
gen_input_real[573] = -32'sd3705;
gen_input_real[829] = -32'sd4765;
gen_input_real[125] = 32'sd2613;
gen_input_real[381] = 32'sd4507;
gen_input_real[637] = 32'sd4217;
gen_input_real[893] = -32'sd5225;
gen_input_real[189] = -32'sd9553;
gen_input_real[445] = 32'sd5631;
gen_input_real[701] = 32'sd8637;
gen_input_real[957] = -32'sd5214;
gen_input_real[253] = -32'sd3868;
gen_input_real[509] = 32'sd5129;
gen_input_real[765] = -32'sd982;
gen_input_real[1021] = -32'sd4183;
gen_input_real[2] = 32'sd4183;
gen_input_real[258] = 32'sd982;
gen_input_real[514] = -32'sd5129;
gen_input_real[770] = 32'sd3868;
gen_input_real[66] = 32'sd5214;
gen_input_real[322] = -32'sd8637;
gen_input_real[578] = -32'sd5631;
gen_input_real[834] = 32'sd9553;
gen_input_real[130] = 32'sd5225;
gen_input_real[386] = -32'sd4217;
gen_input_real[642] = -32'sd4507;
gen_input_real[898] = -32'sd2613;
gen_input_real[194] = 32'sd4765;
gen_input_real[450] = 32'sd3705;
gen_input_real[706] = -32'sd4282;
gen_input_real[962] = -32'sd70;
gen_input_real[18] = 32'sd1394;
gen_input_real[274] = -32'sd1732;
gen_input_real[530] = 32'sd2681;
gen_input_real[786] = 32'sd681;
gen_input_real[82] = -32'sd5434;
gen_input_real[338] = -32'sd149;
gen_input_real[594] = 32'sd4880;
gen_input_real[850] = 32'sd719;
gen_input_real[146] = -32'sd2277;
gen_input_real[402] = -32'sd1588;
gen_input_real[658] = 32'sd2514;
gen_input_real[914] = 32'sd3002;
gen_input_real[210] = -32'sd7510;
gen_input_real[466] = -32'sd3103;
gen_input_real[722] = 32'sd13595;
gen_input_real[978] = -32'sd429;
gen_input_real[34] = -32'sd16704;
gen_input_real[290] = 32'sd5078;
gen_input_real[546] = 32'sd15504;
gen_input_real[802] = -32'sd5778;
gen_input_real[98] = -32'sd10861;
gen_input_real[354] = 32'sd1277;
gen_input_real[610] = 32'sd4727;
gen_input_real[866] = 32'sd3845;
gen_input_real[162] = 32'sd302;
gen_input_real[418] = -32'sd4434;
gen_input_real[674] = -32'sd2587;
gen_input_real[930] = -32'sd241;
gen_input_real[226] = 32'sd2811;
gen_input_real[482] = 32'sd7226;
gen_input_real[738] = -32'sd1795;
gen_input_real[994] = -32'sd10877;
gen_input_real[50] = -32'sd660;
gen_input_real[306] = 32'sd7591;
gen_input_real[562] = 32'sd4066;
gen_input_real[818] = -32'sd2587;
gen_input_real[114] = -32'sd6603;
gen_input_real[370] = 32'sd3311;
gen_input_real[626] = 32'sd6371;
gen_input_real[882] = -32'sd6929;
gen_input_real[178] = -32'sd3176;
gen_input_real[434] = 32'sd5354;
gen_input_real[690] = -32'sd227;
gen_input_real[946] = 32'sd1411;
gen_input_real[242] = 32'sd265;
gen_input_real[498] = -32'sd6368;
gen_input_real[754] = 32'sd3262;
gen_input_real[1010] = 32'sd5970;
gen_input_real[6] = -32'sd7173;
gen_input_real[262] = -32'sd4306;
gen_input_real[518] = 32'sd8711;
gen_input_real[774] = 32'sd6042;
gen_input_real[70] = -32'sd8817;
gen_input_real[326] = -32'sd9930;
gen_input_real[582] = 32'sd9660;
gen_input_real[838] = 32'sd12207;
gen_input_real[134] = -32'sd10422;
gen_input_real[390] = -32'sd10842;
gen_input_real[646] = 32'sd10288;
gen_input_real[902] = 32'sd6215;
gen_input_real[198] = -32'sd8996;
gen_input_real[454] = -32'sd1121;
gen_input_real[710] = 32'sd5215;
gen_input_real[966] = -32'sd426;
gen_input_real[22] = -32'sd1857;
gen_input_real[278] = -32'sd2598;
gen_input_real[534] = 32'sd4054;
gen_input_real[790] = 32'sd5306;
gen_input_real[86] = -32'sd9640;
gen_input_real[342] = -32'sd3127;
gen_input_real[598] = 32'sd12889;
gen_input_real[854] = -32'sd2197;
gen_input_real[150] = -32'sd13843;
gen_input_real[406] = 32'sd6847;
gen_input_real[662] = 32'sd14398;
gen_input_real[918] = -32'sd8031;
gen_input_real[214] = -32'sd13683;
gen_input_real[470] = 32'sd3452;
gen_input_real[726] = 32'sd12329;
gen_input_real[982] = 32'sd4009;
gen_input_real[38] = -32'sd11519;
gen_input_real[294] = -32'sd6881;
gen_input_real[550] = 32'sd8442;
gen_input_real[806] = 32'sd4134;
gen_input_real[102] = -32'sd2061;
gen_input_real[358] = -32'sd2516;
gen_input_real[614] = -32'sd1760;
gen_input_real[870] = 32'sd5892;
gen_input_real[166] = -32'sd154;
gen_input_real[422] = -32'sd10321;
gen_input_real[678] = 32'sd3112;
gen_input_real[934] = 32'sd10514;
gen_input_real[230] = -32'sd4196;
gen_input_real[486] = -32'sd8096;
gen_input_real[742] = 32'sd5086;
gen_input_real[998] = 32'sd8295;
gen_input_real[54] = -32'sd5475;
gen_input_real[310] = -32'sd10664;
gen_input_real[566] = 32'sd3316;
gen_input_real[822] = 32'sd10763;
gen_input_real[118] = 32'sd348;
gen_input_real[374] = -32'sd8644;
gen_input_real[630] = -32'sd2300;
gen_input_real[886] = 32'sd7445;
gen_input_real[182] = 32'sd779;
gen_input_real[438] = -32'sd7378;
gen_input_real[694] = 32'sd4589;
gen_input_real[950] = 32'sd8082;
gen_input_real[246] = -32'sd12818;
gen_input_real[502] = -32'sd10307;
gen_input_real[758] = 32'sd19850;
gen_input_real[1014] = 32'sd12465;
gen_input_real[10] = -32'sd20760;
gen_input_real[266] = -32'sd12351;
gen_input_real[522] = 32'sd15919;
gen_input_real[778] = 32'sd11722;
gen_input_real[74] = -32'sd10409;
gen_input_real[330] = -32'sd12634;
gen_input_real[586] = 32'sd6690;
gen_input_real[842] = 32'sd12151;
gen_input_real[138] = -32'sd5051;
gen_input_real[394] = -32'sd8816;
gen_input_real[650] = 32'sd5754;
gen_input_real[906] = 32'sd6940;
gen_input_real[202] = -32'sd5795;
gen_input_real[458] = -32'sd7787;
gen_input_real[714] = 32'sd2492;
gen_input_real[970] = 32'sd7792;
gen_input_real[26] = 32'sd1076;
gen_input_real[282] = -32'sd7117;
gen_input_real[538] = -32'sd750;
gen_input_real[794] = 32'sd8654;
gen_input_real[90] = -32'sd2563;
gen_input_real[346] = -32'sd9741;
gen_input_real[602] = 32'sd4164;
gen_input_real[858] = 32'sd5576;
gen_input_real[154] = -32'sd1131;
gen_input_real[410] = -32'sd68;
gen_input_real[666] = -32'sd3979;
gen_input_real[922] = 32'sd1106;
gen_input_real[218] = 32'sd6057;
gen_input_real[474] = -32'sd7144;
gen_input_real[730] = -32'sd3518;
gen_input_real[986] = 32'sd12156;
gen_input_real[42] = -32'sd180;
gen_input_real[298] = -32'sd15824;
gen_input_real[554] = 32'sd1590;
gen_input_real[810] = 32'sd17782;
gen_input_real[106] = -32'sd1907;
gen_input_real[362] = -32'sd16626;
gen_input_real[618] = 32'sd3158;
gen_input_real[874] = 32'sd16197;
gen_input_real[170] = -32'sd4268;
gen_input_real[426] = -32'sd19013;
gen_input_real[682] = 32'sd3545;
gen_input_real[938] = 32'sd21128;
gen_input_real[234] = -32'sd413;
gen_input_real[490] = -32'sd19885;
gen_input_real[746] = -32'sd3406;
gen_input_real[1002] = 32'sd17243;
gen_input_real[58] = 32'sd5189;
gen_input_real[314] = -32'sd13938;
gen_input_real[570] = -32'sd5177;
gen_input_real[826] = 32'sd9533;
gen_input_real[122] = 32'sd4027;
gen_input_real[378] = -32'sd7084;
gen_input_real[634] = -32'sd663;
gen_input_real[890] = 32'sd8507;
gen_input_real[186] = -32'sd3926;
gen_input_real[442] = -32'sd10388;
gen_input_real[698] = 32'sd6724;
gen_input_real[954] = 32'sd9833;
gen_input_real[250] = -32'sd6111;
gen_input_real[506] = -32'sd7263;
gen_input_real[762] = 32'sd2703;
gen_input_real[1018] = 32'sd4090;
gen_input_real[14] = 32'sd1168;
gen_input_real[270] = -32'sd2481;
gen_input_real[526] = -32'sd3450;
gen_input_real[782] = 32'sd3393;
gen_input_real[78] = 32'sd4823;
gen_input_real[334] = -32'sd4922;
gen_input_real[590] = -32'sd6110;
gen_input_real[846] = 32'sd6284;
gen_input_real[142] = 32'sd5502;
gen_input_real[398] = -32'sd9381;
gen_input_real[654] = -32'sd3031;
gen_input_real[910] = 32'sd14123;
gen_input_real[206] = 32'sd3026;
gen_input_real[462] = -32'sd17185;
gen_input_real[718] = -32'sd7631;
gen_input_real[974] = 32'sd16411;
gen_input_real[30] = 32'sd13351;
gen_input_real[286] = -32'sd12692;
gen_input_real[542] = -32'sd16277;
gen_input_real[798] = 32'sd7917;
gen_input_real[94] = 32'sd15841;
gen_input_real[350] = -32'sd4349;
gen_input_real[606] = -32'sd13625;
gen_input_real[862] = 32'sd4796;
gen_input_real[158] = 32'sd11315;
gen_input_real[414] = -32'sd9103;
gen_input_real[670] = -32'sd9183;
gen_input_real[926] = 32'sd12171;
gen_input_real[222] = 32'sd6056;
gen_input_real[478] = -32'sd11130;
gen_input_real[734] = -32'sd2447;
gen_input_real[990] = 32'sd9964;
gen_input_real[46] = 32'sd1298;
gen_input_real[302] = -32'sd10997;
gen_input_real[558] = -32'sd2052;
gen_input_real[814] = 32'sd11506;
gen_input_real[110] = 32'sd541;
gen_input_real[366] = -32'sd10478;
gen_input_real[622] = 32'sd2647;
gen_input_real[878] = 32'sd8346;
gen_input_real[174] = -32'sd2372;
gen_input_real[430] = -32'sd4970;
gen_input_real[686] = -32'sd2614;
gen_input_real[942] = 32'sd2648;
gen_input_real[238] = 32'sd7551;
gen_input_real[494] = -32'sd4560;
gen_input_real[750] = -32'sd8701;
gen_input_real[1006] = 32'sd9104;
gen_input_real[62] = 32'sd7780;
gen_input_real[318] = -32'sd10377;
gen_input_real[574] = -32'sd6400;
gen_input_real[830] = 32'sd6063;
gen_input_real[126] = 32'sd5057;
gen_input_real[382] = -32'sd24;
gen_input_real[638] = -32'sd6816;
gen_input_real[894] = -32'sd3789;
gen_input_real[190] = 32'sd11391;
gen_input_real[446] = 32'sd4169;
gen_input_real[702] = -32'sd14342;
gen_input_real[958] = -32'sd2393;
gen_input_real[254] = 32'sd15184;
gen_input_real[510] = 32'sd1638;
gen_input_real[766] = -32'sd14521;
gen_input_real[1022] = -32'sd3307;
gen_input_real[3] = 32'sd10345;
gen_input_real[259] = 32'sd5401;
gen_input_real[515] = -32'sd5154;
gen_input_real[771] = -32'sd3342;
gen_input_real[67] = 32'sd5132;
gen_input_real[323] = -32'sd5404;
gen_input_real[579] = -32'sd8783;
gen_input_real[835] = 32'sd14576;
gen_input_real[131] = 32'sd8588;
gen_input_real[387] = -32'sd15888;
gen_input_real[643] = -32'sd5084;
gen_input_real[899] = 32'sd10570;
gen_input_real[195] = 32'sd5033;
gen_input_real[451] = -32'sd4813;
gen_input_real[707] = -32'sd8309;
gen_input_real[963] = 32'sd1513;
gen_input_real[19] = 32'sd10516;
gen_input_real[275] = -32'sd1376;
gen_input_real[531] = -32'sd10566;
gen_input_real[787] = 32'sd4273;
gen_input_real[83] = 32'sd8386;
gen_input_real[339] = -32'sd7670;
gen_input_real[595] = -32'sd4419;
gen_input_real[851] = 32'sd8111;
gen_input_real[147] = 32'sd1559;
gen_input_real[403] = -32'sd5087;
gen_input_real[659] = -32'sd2009;
gen_input_real[915] = 32'sd705;
gen_input_real[211] = 32'sd4254;
gen_input_real[467] = 32'sd3460;
gen_input_real[723] = -32'sd5029;
gen_input_real[979] = -32'sd6916;
gen_input_real[35] = 32'sd3137;
gen_input_real[291] = 32'sd9462;
gen_input_real[547] = 32'sd250;
gen_input_real[803] = -32'sd10564;
gen_input_real[99] = -32'sd3339;
gen_input_real[355] = 32'sd9484;
gen_input_real[611] = 32'sd3625;
gen_input_real[867] = -32'sd5975;
gen_input_real[163] = 32'sd616;
gen_input_real[419] = 32'sd599;
gen_input_real[675] = -32'sd6513;
gen_input_real[931] = 32'sd3888;
gen_input_real[227] = 32'sd8270;
gen_input_real[483] = -32'sd3840;
gen_input_real[739] = -32'sd5575;
gen_input_real[995] = 32'sd147;
gen_input_real[51] = 32'sd4325;
gen_input_real[307] = 32'sd1951;
gen_input_real[563] = -32'sd7159;
gen_input_real[819] = -32'sd581;
gen_input_real[115] = 32'sd10763;
gen_input_real[371] = 32'sd52;
gen_input_real[627] = -32'sd11599;
gen_input_real[883] = -32'sd2515;
gen_input_real[179] = 32'sd10120;
gen_input_real[435] = 32'sd3785;
gen_input_real[691] = -32'sd9289;
gen_input_real[947] = -32'sd1438;
gen_input_real[243] = 32'sd9058;
gen_input_real[499] = -32'sd1911;
gen_input_real[755] = -32'sd7133;
gen_input_real[1011] = 32'sd3762;
gen_input_real[7] = 32'sd3505;
gen_input_real[263] = -32'sd4242;
gen_input_real[519] = 32'sd1032;
gen_input_real[775] = 32'sd3851;
gen_input_real[71] = -32'sd5372;
gen_input_real[327] = -32'sd1420;
gen_input_real[583] = 32'sd6785;
gen_input_real[839] = -32'sd1881;
gen_input_real[135] = -32'sd4436;
gen_input_real[391] = 32'sd1961;
gen_input_real[647] = 32'sd2152;
gen_input_real[903] = 32'sd496;
gen_input_real[199] = -32'sd3668;
gen_input_real[455] = -32'sd2012;
gen_input_real[711] = 32'sd6701;
gen_input_real[967] = 32'sd3099;
gen_input_real[23] = -32'sd7072;
gen_input_real[279] = -32'sd4006;
gen_input_real[535] = 32'sd4644;
gen_input_real[791] = 32'sd3536;
gen_input_real[87] = 32'sd28;
gen_input_real[343] = -32'sd3136;
gen_input_real[599] = -32'sd5298;
gen_input_real[855] = 32'sd2751;
gen_input_real[151] = 32'sd5951;
gen_input_real[407] = 32'sd1893;
gen_input_real[663] = -32'sd1651;
gen_input_real[919] = -32'sd10997;
gen_input_real[215] = -32'sd1569;
gen_input_real[471] = 32'sd16020;
gen_input_real[727] = 32'sd669;
gen_input_real[983] = -32'sd11455;
gen_input_real[39] = 32'sd2460;
gen_input_real[295] = 32'sd3450;
gen_input_real[551] = -32'sd4464;
gen_input_real[807] = 32'sd1286;
gen_input_real[103] = 32'sd3836;
gen_input_real[359] = -32'sd3143;
gen_input_real[615] = -32'sd1987;
gen_input_real[871] = 32'sd4152;
gen_input_real[167] = 32'sd717;
gen_input_real[423] = -32'sd4643;
gen_input_real[679] = -32'sd280;
gen_input_real[935] = 32'sd3880;
gen_input_real[231] = -32'sd365;
gen_input_real[487] = -32'sd2686;
gen_input_real[743] = 32'sd1567;
gen_input_real[999] = 32'sd3726;
gen_input_real[55] = -32'sd2524;
gen_input_real[311] = -32'sd7464;
gen_input_real[567] = 32'sd2428;
gen_input_real[823] = 32'sd11649;
gen_input_real[119] = -32'sd441;
gen_input_real[375] = -32'sd14036;
gen_input_real[631] = -32'sd2799;
gen_input_real[887] = 32'sd13175;
gen_input_real[183] = 32'sd4542;
gen_input_real[439] = -32'sd9327;
gen_input_real[695] = -32'sd3195;
gen_input_real[951] = 32'sd5455;
gen_input_real[247] = 32'sd73;
gen_input_real[503] = -32'sd3763;
gen_input_real[759] = 32'sd3027;
gen_input_real[1015] = 32'sd2792;
gen_input_real[11] = -32'sd5986;
gen_input_real[267] = -32'sd1033;
gen_input_real[523] = 32'sd8652;
gen_input_real[779] = -32'sd858;
gen_input_real[75] = -32'sd9012;
gen_input_real[331] = 32'sd2814;
gen_input_real[587] = 32'sd6068;
gen_input_real[843] = -32'sd4373;
gen_input_real[139] = -32'sd2464;
gen_input_real[395] = 32'sd2290;
gen_input_real[651] = 32'sd1112;
gen_input_real[907] = 32'sd4739;
gen_input_real[203] = -32'sd1788;
gen_input_real[459] = -32'sd11210;
gen_input_real[715] = 32'sd2637;
gen_input_real[971] = 32'sd10150;
gen_input_real[27] = -32'sd2278;
gen_input_real[283] = -32'sd3719;
gen_input_real[539] = -32'sd550;
gen_input_real[795] = 32'sd856;
gen_input_real[91] = 32'sd5202;
gen_input_real[347] = -32'sd3608;
gen_input_real[603] = -32'sd7577;
gen_input_real[859] = 32'sd6889;
gen_input_real[155] = 32'sd6885;
gen_input_real[411] = -32'sd7734;
gen_input_real[667] = -32'sd6876;
gen_input_real[923] = 32'sd6765;
gen_input_real[219] = 32'sd8256;
gen_input_real[475] = -32'sd6405;
gen_input_real[731] = -32'sd9584;
gen_input_real[987] = 32'sd8743;
gen_input_real[43] = 32'sd10300;
gen_input_real[299] = -32'sd12457;
gen_input_real[555] = -32'sd9790;
gen_input_real[811] = 32'sd12626;
gen_input_real[107] = 32'sd7160;
gen_input_real[363] = -32'sd7784;
gen_input_real[619] = -32'sd1392;
gen_input_real[875] = 32'sd4135;
gen_input_real[171] = -32'sd5422;
gen_input_real[427] = -32'sd4955;
gen_input_real[683] = 32'sd8371;
gen_input_real[939] = 32'sd7124;
gen_input_real[235] = -32'sd6270;
gen_input_real[491] = -32'sd10472;
gen_input_real[747] = 32'sd2287;
gen_input_real[1003] = 32'sd15024;
gen_input_real[59] = 32'sd1237;
gen_input_real[315] = -32'sd16469;
gen_input_real[571] = -32'sd4207;
gen_input_real[827] = 32'sd13848;
gen_input_real[123] = 32'sd5640;
gen_input_real[379] = -32'sd10494;
gen_input_real[635] = -32'sd3798;
gen_input_real[891] = 32'sd7539;
gen_input_real[187] = 32'sd863;
gen_input_real[443] = -32'sd4581;
gen_input_real[699] = -32'sd696;
gen_input_real[955] = 32'sd2373;
gen_input_real[251] = 32'sd3003;
gen_input_real[507] = -32'sd1521;
gen_input_real[763] = -32'sd6293;
gen_input_real[1019] = 32'sd1261;
gen_input_real[15] = 32'sd9697;
gen_input_real[271] = -32'sd1478;
gen_input_real[527] = -32'sd11372;
gen_input_real[783] = 32'sd2298;
gen_input_real[79] = 32'sd12016;
gen_input_real[335] = -32'sd1544;
gen_input_real[591] = -32'sd13369;
gen_input_real[847] = -32'sd552;
gen_input_real[143] = 32'sd13556;
gen_input_real[399] = -32'sd355;
gen_input_real[655] = -32'sd9956;
gen_input_real[911] = 32'sd5124;
gen_input_real[207] = 32'sd4224;
gen_input_real[463] = -32'sd9279;
gen_input_real[719] = -32'sd1896;
gen_input_real[975] = 32'sd9771;
gen_input_real[31] = 32'sd5676;
gen_input_real[287] = -32'sd9027;
gen_input_real[543] = -32'sd11486;
gen_input_real[799] = 32'sd9909;
gen_input_real[95] = 32'sd13410;
gen_input_real[351] = -32'sd11578;
gen_input_real[607] = -32'sd11736;
gen_input_real[863] = 32'sd12980;
gen_input_real[159] = 32'sd12014;
gen_input_real[415] = -32'sd13828;
gen_input_real[671] = -32'sd14897;
gen_input_real[927] = 32'sd13278;
gen_input_real[223] = 32'sd15447;
gen_input_real[479] = -32'sd11291;
gen_input_real[735] = -32'sd11915;
gen_input_real[991] = 32'sd8610;
gen_input_real[47] = 32'sd7215;
gen_input_real[303] = -32'sd4629;
gen_input_real[559] = -32'sd3916;
gen_input_real[815] = -32'sd841;
gen_input_real[111] = 32'sd2677;
gen_input_real[367] = 32'sd4015;
gen_input_real[623] = -32'sd4429;
gen_input_real[879] = -32'sd2125;
gen_input_real[175] = 32'sd8359;
gen_input_real[431] = -32'sd1536;
gen_input_real[687] = -32'sd9639;
gen_input_real[943] = 32'sd2951;
gen_input_real[239] = 32'sd6746;
gen_input_real[495] = -32'sd1236;
gen_input_real[751] = -32'sd5221;
gen_input_real[1007] = -32'sd2436;
gen_input_real[63] = 32'sd7812;
gen_input_real[319] = 32'sd4364;
gen_input_real[575] = -32'sd10567;
gen_input_real[831] = -32'sd2032;
gen_input_real[127] = 32'sd10725;
gen_input_real[383] = -32'sd2057;
gen_input_real[639] = -32'sd9073;
gen_input_real[895] = 32'sd4174;
gen_input_real[191] = 32'sd7035;
gen_input_real[447] = -32'sd2547;
gen_input_real[703] = -32'sd8653;
gen_input_real[959] = -32'sd963;
gen_input_real[255] = 32'sd19335;
gen_input_real[511] = 32'sd2085;
gen_input_real[767] = -32'sd32767;
gen_input_real[1023] = 32'sd0;
