gen_input_real[0] = 16'sd0;
gen_input_real[16] = 16'sd127;
gen_input_real[32] = -16'sd26;
gen_input_real[48] = -16'sd94;
gen_input_real[4] = 16'sd37;
gen_input_real[20] = 16'sd58;
gen_input_real[36] = -16'sd39;
gen_input_real[52] = -16'sd30;
gen_input_real[8] = 16'sd41;
gen_input_real[24] = 16'sd13;
gen_input_real[40] = -16'sd45;
gen_input_real[56] = -16'sd7;
gen_input_real[12] = 16'sd42;
gen_input_real[28] = 16'sd3;
gen_input_real[44] = -16'sd28;
gen_input_real[60] = -16'sd5;
gen_input_real[1] = 16'sd8;
gen_input_real[17] = 16'sd9;
gen_input_real[33] = 16'sd9;
gen_input_real[49] = -16'sd7;
gen_input_real[5] = -16'sd17;
gen_input_real[21] = -16'sd2;
gen_input_real[37] = 16'sd16;
gen_input_real[53] = 16'sd16;
gen_input_real[9] = -16'sd14;
gen_input_real[25] = -16'sd25;
gen_input_real[41] = 16'sd13;
gen_input_real[57] = 16'sd17;
gen_input_real[13] = -16'sd8;
gen_input_real[29] = 16'sd2;
gen_input_real[45] = -16'sd3;
gen_input_real[61] = -16'sd11;
gen_input_real[2] = 16'sd11;
gen_input_real[18] = 16'sd3;
gen_input_real[34] = -16'sd2;
gen_input_real[50] = 16'sd8;
gen_input_real[6] = -16'sd17;
gen_input_real[22] = -16'sd13;
gen_input_real[38] = 16'sd25;
gen_input_real[54] = 16'sd14;
gen_input_real[10] = -16'sd16;
gen_input_real[26] = -16'sd16;
gen_input_real[42] = 16'sd2;
gen_input_real[58] = 16'sd17;
gen_input_real[14] = 16'sd7;
gen_input_real[30] = -16'sd9;
gen_input_real[46] = -16'sd9;
gen_input_real[62] = -16'sd8;
gen_input_real[3] = 16'sd5;
gen_input_real[19] = 16'sd28;
gen_input_real[35] = -16'sd3;
gen_input_real[51] = -16'sd42;
gen_input_real[7] = 16'sd7;
gen_input_real[23] = 16'sd45;
gen_input_real[39] = -16'sd13;
gen_input_real[55] = -16'sd41;
gen_input_real[11] = 16'sd30;
gen_input_real[27] = 16'sd39;
gen_input_real[43] = -16'sd58;
gen_input_real[59] = -16'sd37;
gen_input_real[15] = 16'sd94;
gen_input_real[31] = 16'sd26;
gen_input_real[47] = -16'sd127;
gen_input_real[63] = 16'sd0;
