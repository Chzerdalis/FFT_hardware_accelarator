0 0
10 -54
68 -164
234 -351
912 -912
-366 245
-342 141
-354 70
-324 0
-354 -70
-342 -141
-366 -245
912 912
234 351
68 164
10 54
