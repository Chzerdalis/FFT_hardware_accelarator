0 0
4 -99
20 -204
51 -350
99 -502
201 -805
188 -620
283 -792
404 -975
576 -1219
835 -1563
1325 -2212
4689 -7019
752 -1014
2263 -2758
7822 -8631
8118 -8118
9517 -8626
3152 -2587
-3240 2403
-3111 2079
-4578 2744
-1416 757
-4439 2099
-2970 1230
-3326 1190
-2778 842
-2772 694
-2654 527
-2682 397
-2560 252
-2522 123
-2512 0
-2522 -123
-2560 -252
-2682 -397
-2654 -527
-2772 -694
-2778 -842
-3326 -1190
-2970 -1230
-4439 -2099
-1416 -757
-4578 -2744
-3111 -2079
-3240 -2403
3152 2587
9517 8626
8118 8118
7822 8631
2263 2758
752 1014
4689 7019
1325 2212
835 1563
576 1219
404 975
283 792
188 620
201 805
99 502
51 350
20 204
4 99
