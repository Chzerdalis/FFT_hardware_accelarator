gen_input_real[0] = 24'sd0;
gen_input_real[64] = 24'sd2047;
gen_input_real[128] = -24'sd38;
gen_input_real[192] = -24'sd1625;
gen_input_real[16] = 24'sd99;
gen_input_real[80] = 24'sd1218;
gen_input_real[144] = -24'sd170;
gen_input_real[208] = -24'sd995;
gen_input_real[32] = 24'sd244;
gen_input_real[96] = 24'sd813;
gen_input_real[160] = -24'sd353;
gen_input_real[224] = -24'sd571;
gen_input_real[48] = 24'sd490;
gen_input_real[112] = 24'sd385;
gen_input_real[176] = -24'sd593;
gen_input_real[240] = -24'sd442;
gen_input_real[4] = 24'sd592;
gen_input_real[68] = 24'sd645;
gen_input_real[132] = -24'sd511;
gen_input_real[196] = -24'sd708;
gen_input_real[20] = 24'sd499;
gen_input_real[84] = 24'sd498;
gen_input_real[148] = -24'sd579;
gen_input_real[212] = -24'sd107;
gen_input_real[36] = 24'sd620;
gen_input_real[100] = -24'sd248;
gen_input_real[164] = -24'sd614;
gen_input_real[228] = 24'sd500;
gen_input_real[52] = 24'sd637;
gen_input_real[116] = -24'sd730;
gen_input_real[180] = -24'sd692;
gen_input_real[244] = 24'sd900;
gen_input_real[8] = 24'sd748;
gen_input_real[72] = -24'sd874;
gen_input_real[136] = -24'sd760;
gen_input_real[200] = 24'sd619;
gen_input_real[24] = 24'sd692;
gen_input_real[88] = -24'sd300;
gen_input_real[152] = -24'sd565;
gen_input_real[216] = 24'sd116;
gen_input_real[40] = 24'sd492;
gen_input_real[104] = -24'sd59;
gen_input_real[168] = -24'sd554;
gen_input_real[232] = 24'sd61;
gen_input_real[56] = 24'sd626;
gen_input_real[120] = -24'sd134;
gen_input_real[184] = -24'sd599;
gen_input_real[248] = 24'sd273;
gen_input_real[12] = 24'sd546;
gen_input_real[76] = -24'sd424;
gen_input_real[140] = -24'sd537;
gen_input_real[204] = 24'sd466;
gen_input_real[28] = 24'sd529;
gen_input_real[92] = -24'sd318;
gen_input_real[156] = -24'sd424;
gen_input_real[220] = 24'sd105;
gen_input_real[44] = 24'sd239;
gen_input_real[108] = 24'sd23;
gen_input_real[172] = -24'sd104;
gen_input_real[236] = -24'sd125;
gen_input_real[60] = 24'sd40;
gen_input_real[124] = 24'sd252;
gen_input_real[188] = -24'sd21;
gen_input_real[252] = -24'sd278;
gen_input_real[1] = 24'sd54;
gen_input_real[65] = 24'sd120;
gen_input_real[129] = -24'sd74;
gen_input_real[193] = 24'sd113;
gen_input_real[17] = 24'sd36;
gen_input_real[81] = -24'sd276;
gen_input_real[145] = 24'sd23;
gen_input_real[209] = 24'sd347;
gen_input_real[33] = -24'sd109;
gen_input_real[97] = -24'sd371;
gen_input_real[161] = 24'sd217;
gen_input_real[225] = 24'sd340;
gen_input_real[49] = -24'sd307;
gen_input_real[113] = -24'sd240;
gen_input_real[177] = 24'sd359;
gen_input_real[241] = 24'sd133;
gen_input_real[5] = -24'sd337;
gen_input_real[69] = -24'sd49;
gen_input_real[133] = 24'sd214;
gen_input_real[197] = -24'sd21;
gen_input_real[21] = -24'sd33;
gen_input_real[85] = 24'sd31;
gen_input_real[149] = -24'sd125;
gen_input_real[213] = 24'sd67;
gen_input_real[37] = 24'sd228;
gen_input_real[101] = -24'sd205;
gen_input_real[165] = -24'sd285;
gen_input_real[229] = 24'sd302;
gen_input_real[53] = 24'sd271;
gen_input_real[117] = -24'sd351;
gen_input_real[181] = -24'sd187;
gen_input_real[245] = 24'sd350;
gen_input_real[9] = 24'sd135;
gen_input_real[73] = -24'sd300;
gen_input_real[137] = -24'sd183;
gen_input_real[201] = 24'sd262;
gen_input_real[25] = 24'sd275;
gen_input_real[89] = -24'sd245;
gen_input_real[153] = -24'sd342;
gen_input_real[217] = 24'sd186;
gen_input_real[41] = 24'sd422;
gen_input_real[105] = -24'sd125;
gen_input_real[169] = -24'sd548;
gen_input_real[233] = 24'sd184;
gen_input_real[57] = 24'sd623;
gen_input_real[121] = -24'sd390;
gen_input_real[185] = -24'sd522;
gen_input_real[249] = 24'sd630;
gen_input_real[13] = 24'sd290;
gen_input_real[77] = -24'sd751;
gen_input_real[141] = -24'sd45;
gen_input_real[205] = 24'sd751;
gen_input_real[29] = -24'sd154;
gen_input_real[93] = -24'sd758;
gen_input_real[157] = 24'sd259;
gen_input_real[221] = 24'sd806;
gen_input_real[45] = -24'sd296;
gen_input_real[109] = -24'sd763;
gen_input_real[173] = 24'sd369;
gen_input_real[237] = 24'sd550;
gen_input_real[61] = -24'sd430;
gen_input_real[125] = -24'sd317;
gen_input_real[189] = 24'sd365;
gen_input_real[253] = 24'sd261;
gen_input_real[2] = -24'sd261;
gen_input_real[66] = -24'sd365;
gen_input_real[130] = 24'sd317;
gen_input_real[194] = 24'sd430;
gen_input_real[18] = -24'sd550;
gen_input_real[82] = -24'sd369;
gen_input_real[146] = 24'sd763;
gen_input_real[210] = 24'sd296;
gen_input_real[34] = -24'sd806;
gen_input_real[98] = -24'sd259;
gen_input_real[162] = 24'sd758;
gen_input_real[226] = 24'sd154;
gen_input_real[50] = -24'sd751;
gen_input_real[114] = 24'sd45;
gen_input_real[178] = 24'sd751;
gen_input_real[242] = -24'sd290;
gen_input_real[6] = -24'sd630;
gen_input_real[70] = 24'sd522;
gen_input_real[134] = 24'sd390;
gen_input_real[198] = -24'sd623;
gen_input_real[22] = -24'sd184;
gen_input_real[86] = 24'sd548;
gen_input_real[150] = 24'sd125;
gen_input_real[214] = -24'sd422;
gen_input_real[38] = -24'sd186;
gen_input_real[102] = 24'sd342;
gen_input_real[166] = 24'sd245;
gen_input_real[230] = -24'sd275;
gen_input_real[54] = -24'sd262;
gen_input_real[118] = 24'sd183;
gen_input_real[182] = 24'sd300;
gen_input_real[246] = -24'sd135;
gen_input_real[10] = -24'sd350;
gen_input_real[74] = 24'sd187;
gen_input_real[138] = 24'sd351;
gen_input_real[202] = -24'sd271;
gen_input_real[26] = -24'sd302;
gen_input_real[90] = 24'sd285;
gen_input_real[154] = 24'sd205;
gen_input_real[218] = -24'sd228;
gen_input_real[42] = -24'sd67;
gen_input_real[106] = 24'sd125;
gen_input_real[170] = -24'sd31;
gen_input_real[234] = 24'sd33;
gen_input_real[58] = 24'sd21;
gen_input_real[122] = -24'sd214;
gen_input_real[186] = 24'sd49;
gen_input_real[250] = 24'sd337;
gen_input_real[14] = -24'sd133;
gen_input_real[78] = -24'sd359;
gen_input_real[142] = 24'sd240;
gen_input_real[206] = 24'sd307;
gen_input_real[30] = -24'sd340;
gen_input_real[94] = -24'sd217;
gen_input_real[158] = 24'sd371;
gen_input_real[222] = 24'sd109;
gen_input_real[46] = -24'sd347;
gen_input_real[110] = -24'sd23;
gen_input_real[174] = 24'sd276;
gen_input_real[238] = -24'sd36;
gen_input_real[62] = -24'sd113;
gen_input_real[126] = 24'sd74;
gen_input_real[190] = -24'sd120;
gen_input_real[254] = -24'sd54;
gen_input_real[3] = 24'sd278;
gen_input_real[67] = 24'sd21;
gen_input_real[131] = -24'sd252;
gen_input_real[195] = -24'sd40;
gen_input_real[19] = 24'sd125;
gen_input_real[83] = 24'sd104;
gen_input_real[147] = -24'sd23;
gen_input_real[211] = -24'sd239;
gen_input_real[35] = -24'sd105;
gen_input_real[99] = 24'sd424;
gen_input_real[163] = 24'sd318;
gen_input_real[227] = -24'sd529;
gen_input_real[51] = -24'sd466;
gen_input_real[115] = 24'sd537;
gen_input_real[179] = 24'sd424;
gen_input_real[243] = -24'sd546;
gen_input_real[7] = -24'sd273;
gen_input_real[71] = 24'sd599;
gen_input_real[135] = 24'sd134;
gen_input_real[199] = -24'sd626;
gen_input_real[23] = -24'sd61;
gen_input_real[87] = 24'sd554;
gen_input_real[151] = 24'sd59;
gen_input_real[215] = -24'sd492;
gen_input_real[39] = -24'sd116;
gen_input_real[103] = 24'sd565;
gen_input_real[167] = 24'sd300;
gen_input_real[231] = -24'sd692;
gen_input_real[55] = -24'sd619;
gen_input_real[119] = 24'sd760;
gen_input_real[183] = 24'sd874;
gen_input_real[247] = -24'sd748;
gen_input_real[11] = -24'sd900;
gen_input_real[75] = 24'sd692;
gen_input_real[139] = 24'sd730;
gen_input_real[203] = -24'sd637;
gen_input_real[27] = -24'sd500;
gen_input_real[91] = 24'sd614;
gen_input_real[155] = 24'sd248;
gen_input_real[219] = -24'sd620;
gen_input_real[43] = 24'sd107;
gen_input_real[107] = 24'sd579;
gen_input_real[171] = -24'sd498;
gen_input_real[235] = -24'sd499;
gen_input_real[59] = 24'sd708;
gen_input_real[123] = 24'sd511;
gen_input_real[187] = -24'sd645;
gen_input_real[251] = -24'sd592;
gen_input_real[15] = 24'sd442;
gen_input_real[79] = 24'sd593;
gen_input_real[143] = -24'sd385;
gen_input_real[207] = -24'sd490;
gen_input_real[31] = 24'sd571;
gen_input_real[95] = 24'sd353;
gen_input_real[159] = -24'sd813;
gen_input_real[223] = -24'sd244;
gen_input_real[47] = 24'sd995;
gen_input_real[111] = 24'sd170;
gen_input_real[175] = -24'sd1218;
gen_input_real[239] = -24'sd99;
gen_input_real[63] = 24'sd1625;
gen_input_real[127] = 24'sd38;
gen_input_real[191] = -24'sd2047;
gen_input_real[255] = 24'sd0;
