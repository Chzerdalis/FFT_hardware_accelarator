w_real[0] = 8'h7F; w_imag[0] = 8'h00;
w_real[1] = 8'h7F; w_imag[1] = 8'hFD;
w_real[2] = 8'h7F; w_imag[2] = 8'hFA;
w_real[3] = 8'h7F; w_imag[3] = 8'hF7;
w_real[4] = 8'h7F; w_imag[4] = 8'hF4;
w_real[5] = 8'h7F; w_imag[5] = 8'hF1;
w_real[6] = 8'h7E; w_imag[6] = 8'hEE;
w_real[7] = 8'h7E; w_imag[7] = 8'hEB;
w_real[8] = 8'h7D; w_imag[8] = 8'hE8;
w_real[9] = 8'h7C; w_imag[9] = 8'hE4;
w_real[10] = 8'h7C; w_imag[10] = 8'hE1;
w_real[11] = 8'h7B; w_imag[11] = 8'hDE;
w_real[12] = 8'h7A; w_imag[12] = 8'hDB;
w_real[13] = 8'h79; w_imag[13] = 8'hD8;
w_real[14] = 8'h78; w_imag[14] = 8'hD5;
w_real[15] = 8'h77; w_imag[15] = 8'hD2;
w_real[16] = 8'h76; w_imag[16] = 8'hD0;
w_real[17] = 8'h75; w_imag[17] = 8'hCD;
w_real[18] = 8'h73; w_imag[18] = 8'hCA;
w_real[19] = 8'h72; w_imag[19] = 8'hC7;
w_real[20] = 8'h70; w_imag[20] = 8'hC4;
w_real[21] = 8'h6F; w_imag[21] = 8'hC1;
w_real[22] = 8'h6D; w_imag[22] = 8'hBF;
w_real[23] = 8'h6C; w_imag[23] = 8'hBC;
w_real[24] = 8'h6A; w_imag[24] = 8'hB9;
w_real[25] = 8'h68; w_imag[25] = 8'hB7;
w_real[26] = 8'h66; w_imag[26] = 8'hB4;
w_real[27] = 8'h64; w_imag[27] = 8'hB2;
w_real[28] = 8'h62; w_imag[28] = 8'hAF;
w_real[29] = 8'h60; w_imag[29] = 8'hAD;
w_real[30] = 8'h5E; w_imag[30] = 8'hAB;
w_real[31] = 8'h5C; w_imag[31] = 8'hA8;
w_real[32] = 8'h5A; w_imag[32] = 8'hA6;
w_real[33] = 8'h58; w_imag[33] = 8'hA4;
w_real[34] = 8'h55; w_imag[34] = 8'hA2;
w_real[35] = 8'h53; w_imag[35] = 8'hA0;
w_real[36] = 8'h51; w_imag[36] = 8'h9E;
w_real[37] = 8'h4E; w_imag[37] = 8'h9C;
w_real[38] = 8'h4C; w_imag[38] = 8'h9A;
w_real[39] = 8'h49; w_imag[39] = 8'h98;
w_real[40] = 8'h47; w_imag[40] = 8'h96;
w_real[41] = 8'h44; w_imag[41] = 8'h94;
w_real[42] = 8'h41; w_imag[42] = 8'h93;
w_real[43] = 8'h3F; w_imag[43] = 8'h91;
w_real[44] = 8'h3C; w_imag[44] = 8'h90;
w_real[45] = 8'h39; w_imag[45] = 8'h8E;
w_real[46] = 8'h36; w_imag[46] = 8'h8D;
w_real[47] = 8'h33; w_imag[47] = 8'h8B;
w_real[48] = 8'h30; w_imag[48] = 8'h8A;
w_real[49] = 8'h2E; w_imag[49] = 8'h89;
w_real[50] = 8'h2B; w_imag[50] = 8'h88;
w_real[51] = 8'h28; w_imag[51] = 8'h87;
w_real[52] = 8'h25; w_imag[52] = 8'h86;
w_real[53] = 8'h22; w_imag[53] = 8'h85;
w_real[54] = 8'h1F; w_imag[54] = 8'h84;
w_real[55] = 8'h1C; w_imag[55] = 8'h84;
w_real[56] = 8'h18; w_imag[56] = 8'h83;
w_real[57] = 8'h15; w_imag[57] = 8'h82;
w_real[58] = 8'h12; w_imag[58] = 8'h82;
w_real[59] = 8'h0F; w_imag[59] = 8'h81;
w_real[60] = 8'h0C; w_imag[60] = 8'h81;
w_real[61] = 8'h09; w_imag[61] = 8'h81;
w_real[62] = 8'h06; w_imag[62] = 8'h81;
w_real[63] = 8'h03; w_imag[63] = 8'h81;
w_real[64] = 8'h00; w_imag[64] = 8'h80;
w_real[65] = 8'hFD; w_imag[65] = 8'h81;
w_real[66] = 8'hFA; w_imag[66] = 8'h81;
w_real[67] = 8'hF7; w_imag[67] = 8'h81;
w_real[68] = 8'hF4; w_imag[68] = 8'h81;
w_real[69] = 8'hF1; w_imag[69] = 8'h81;
w_real[70] = 8'hEE; w_imag[70] = 8'h82;
w_real[71] = 8'hEB; w_imag[71] = 8'h82;
w_real[72] = 8'hE8; w_imag[72] = 8'h83;
w_real[73] = 8'hE4; w_imag[73] = 8'h84;
w_real[74] = 8'hE1; w_imag[74] = 8'h84;
w_real[75] = 8'hDE; w_imag[75] = 8'h85;
w_real[76] = 8'hDB; w_imag[76] = 8'h86;
w_real[77] = 8'hD8; w_imag[77] = 8'h87;
w_real[78] = 8'hD5; w_imag[78] = 8'h88;
w_real[79] = 8'hD2; w_imag[79] = 8'h89;
w_real[80] = 8'hD0; w_imag[80] = 8'h8A;
w_real[81] = 8'hCD; w_imag[81] = 8'h8B;
w_real[82] = 8'hCA; w_imag[82] = 8'h8D;
w_real[83] = 8'hC7; w_imag[83] = 8'h8E;
w_real[84] = 8'hC4; w_imag[84] = 8'h90;
w_real[85] = 8'hC1; w_imag[85] = 8'h91;
w_real[86] = 8'hBF; w_imag[86] = 8'h93;
w_real[87] = 8'hBC; w_imag[87] = 8'h94;
w_real[88] = 8'hB9; w_imag[88] = 8'h96;
w_real[89] = 8'hB7; w_imag[89] = 8'h98;
w_real[90] = 8'hB4; w_imag[90] = 8'h9A;
w_real[91] = 8'hB2; w_imag[91] = 8'h9C;
w_real[92] = 8'hAF; w_imag[92] = 8'h9E;
w_real[93] = 8'hAD; w_imag[93] = 8'hA0;
w_real[94] = 8'hAB; w_imag[94] = 8'hA2;
w_real[95] = 8'hA8; w_imag[95] = 8'hA4;
w_real[96] = 8'hA6; w_imag[96] = 8'hA6;
w_real[97] = 8'hA4; w_imag[97] = 8'hA8;
w_real[98] = 8'hA2; w_imag[98] = 8'hAB;
w_real[99] = 8'hA0; w_imag[99] = 8'hAD;
w_real[100] = 8'h9E; w_imag[100] = 8'hAF;
w_real[101] = 8'h9C; w_imag[101] = 8'hB2;
w_real[102] = 8'h9A; w_imag[102] = 8'hB4;
w_real[103] = 8'h98; w_imag[103] = 8'hB7;
w_real[104] = 8'h96; w_imag[104] = 8'hB9;
w_real[105] = 8'h94; w_imag[105] = 8'hBC;
w_real[106] = 8'h93; w_imag[106] = 8'hBF;
w_real[107] = 8'h91; w_imag[107] = 8'hC1;
w_real[108] = 8'h90; w_imag[108] = 8'hC4;
w_real[109] = 8'h8E; w_imag[109] = 8'hC7;
w_real[110] = 8'h8D; w_imag[110] = 8'hCA;
w_real[111] = 8'h8B; w_imag[111] = 8'hCD;
w_real[112] = 8'h8A; w_imag[112] = 8'hD0;
w_real[113] = 8'h89; w_imag[113] = 8'hD2;
w_real[114] = 8'h88; w_imag[114] = 8'hD5;
w_real[115] = 8'h87; w_imag[115] = 8'hD8;
w_real[116] = 8'h86; w_imag[116] = 8'hDB;
w_real[117] = 8'h85; w_imag[117] = 8'hDE;
w_real[118] = 8'h84; w_imag[118] = 8'hE1;
w_real[119] = 8'h84; w_imag[119] = 8'hE4;
w_real[120] = 8'h83; w_imag[120] = 8'hE8;
w_real[121] = 8'h82; w_imag[121] = 8'hEB;
w_real[122] = 8'h82; w_imag[122] = 8'hEE;
w_real[123] = 8'h81; w_imag[123] = 8'hF1;
w_real[124] = 8'h81; w_imag[124] = 8'hF4;
w_real[125] = 8'h81; w_imag[125] = 8'hF7;
w_real[126] = 8'h81; w_imag[126] = 8'hFA;
w_real[127] = 8'h81; w_imag[127] = 8'hFD;
w_real[128] = 8'h80; w_imag[128] = 8'h00;
w_real[129] = 8'h81; w_imag[129] = 8'h03;
w_real[130] = 8'h81; w_imag[130] = 8'h06;
w_real[131] = 8'h81; w_imag[131] = 8'h09;
w_real[132] = 8'h81; w_imag[132] = 8'h0C;
w_real[133] = 8'h81; w_imag[133] = 8'h0F;
w_real[134] = 8'h82; w_imag[134] = 8'h12;
w_real[135] = 8'h82; w_imag[135] = 8'h15;
w_real[136] = 8'h83; w_imag[136] = 8'h18;
w_real[137] = 8'h84; w_imag[137] = 8'h1C;
w_real[138] = 8'h84; w_imag[138] = 8'h1F;
w_real[139] = 8'h85; w_imag[139] = 8'h22;
w_real[140] = 8'h86; w_imag[140] = 8'h25;
w_real[141] = 8'h87; w_imag[141] = 8'h28;
w_real[142] = 8'h88; w_imag[142] = 8'h2B;
w_real[143] = 8'h89; w_imag[143] = 8'h2E;
w_real[144] = 8'h8A; w_imag[144] = 8'h30;
w_real[145] = 8'h8B; w_imag[145] = 8'h33;
w_real[146] = 8'h8D; w_imag[146] = 8'h36;
w_real[147] = 8'h8E; w_imag[147] = 8'h39;
w_real[148] = 8'h90; w_imag[148] = 8'h3C;
w_real[149] = 8'h91; w_imag[149] = 8'h3F;
w_real[150] = 8'h93; w_imag[150] = 8'h41;
w_real[151] = 8'h94; w_imag[151] = 8'h44;
w_real[152] = 8'h96; w_imag[152] = 8'h47;
w_real[153] = 8'h98; w_imag[153] = 8'h49;
w_real[154] = 8'h9A; w_imag[154] = 8'h4C;
w_real[155] = 8'h9C; w_imag[155] = 8'h4E;
w_real[156] = 8'h9E; w_imag[156] = 8'h51;
w_real[157] = 8'hA0; w_imag[157] = 8'h53;
w_real[158] = 8'hA2; w_imag[158] = 8'h55;
w_real[159] = 8'hA4; w_imag[159] = 8'h58;
w_real[160] = 8'hA6; w_imag[160] = 8'h5A;
w_real[161] = 8'hA8; w_imag[161] = 8'h5C;
w_real[162] = 8'hAB; w_imag[162] = 8'h5E;
w_real[163] = 8'hAD; w_imag[163] = 8'h60;
w_real[164] = 8'hAF; w_imag[164] = 8'h62;
w_real[165] = 8'hB2; w_imag[165] = 8'h64;
w_real[166] = 8'hB4; w_imag[166] = 8'h66;
w_real[167] = 8'hB7; w_imag[167] = 8'h68;
w_real[168] = 8'hB9; w_imag[168] = 8'h6A;
w_real[169] = 8'hBC; w_imag[169] = 8'h6C;
w_real[170] = 8'hBF; w_imag[170] = 8'h6D;
w_real[171] = 8'hC1; w_imag[171] = 8'h6F;
w_real[172] = 8'hC4; w_imag[172] = 8'h70;
w_real[173] = 8'hC7; w_imag[173] = 8'h72;
w_real[174] = 8'hCA; w_imag[174] = 8'h73;
w_real[175] = 8'hCD; w_imag[175] = 8'h75;
w_real[176] = 8'hD0; w_imag[176] = 8'h76;
w_real[177] = 8'hD2; w_imag[177] = 8'h77;
w_real[178] = 8'hD5; w_imag[178] = 8'h78;
w_real[179] = 8'hD8; w_imag[179] = 8'h79;
w_real[180] = 8'hDB; w_imag[180] = 8'h7A;
w_real[181] = 8'hDE; w_imag[181] = 8'h7B;
w_real[182] = 8'hE1; w_imag[182] = 8'h7C;
w_real[183] = 8'hE4; w_imag[183] = 8'h7C;
w_real[184] = 8'hE8; w_imag[184] = 8'h7D;
w_real[185] = 8'hEB; w_imag[185] = 8'h7E;
w_real[186] = 8'hEE; w_imag[186] = 8'h7E;
w_real[187] = 8'hF1; w_imag[187] = 8'h7F;
w_real[188] = 8'hF4; w_imag[188] = 8'h7F;
w_real[189] = 8'hF7; w_imag[189] = 8'h7F;
w_real[190] = 8'hFA; w_imag[190] = 8'h7F;
w_real[191] = 8'hFD; w_imag[191] = 8'h7F;
w_real[192] = 8'h00; w_imag[192] = 8'h7F;
w_real[193] = 8'h03; w_imag[193] = 8'h7F;
w_real[194] = 8'h06; w_imag[194] = 8'h7F;
w_real[195] = 8'h09; w_imag[195] = 8'h7F;
w_real[196] = 8'h0C; w_imag[196] = 8'h7F;
w_real[197] = 8'h0F; w_imag[197] = 8'h7F;
w_real[198] = 8'h12; w_imag[198] = 8'h7E;
w_real[199] = 8'h15; w_imag[199] = 8'h7E;
w_real[200] = 8'h18; w_imag[200] = 8'h7D;
w_real[201] = 8'h1C; w_imag[201] = 8'h7C;
w_real[202] = 8'h1F; w_imag[202] = 8'h7C;
w_real[203] = 8'h22; w_imag[203] = 8'h7B;
w_real[204] = 8'h25; w_imag[204] = 8'h7A;
w_real[205] = 8'h28; w_imag[205] = 8'h79;
w_real[206] = 8'h2B; w_imag[206] = 8'h78;
w_real[207] = 8'h2E; w_imag[207] = 8'h77;
w_real[208] = 8'h30; w_imag[208] = 8'h76;
w_real[209] = 8'h33; w_imag[209] = 8'h75;
w_real[210] = 8'h36; w_imag[210] = 8'h73;
w_real[211] = 8'h39; w_imag[211] = 8'h72;
w_real[212] = 8'h3C; w_imag[212] = 8'h70;
w_real[213] = 8'h3F; w_imag[213] = 8'h6F;
w_real[214] = 8'h41; w_imag[214] = 8'h6D;
w_real[215] = 8'h44; w_imag[215] = 8'h6C;
w_real[216] = 8'h47; w_imag[216] = 8'h6A;
w_real[217] = 8'h49; w_imag[217] = 8'h68;
w_real[218] = 8'h4C; w_imag[218] = 8'h66;
w_real[219] = 8'h4E; w_imag[219] = 8'h64;
w_real[220] = 8'h51; w_imag[220] = 8'h62;
w_real[221] = 8'h53; w_imag[221] = 8'h60;
w_real[222] = 8'h55; w_imag[222] = 8'h5E;
w_real[223] = 8'h58; w_imag[223] = 8'h5C;
w_real[224] = 8'h5A; w_imag[224] = 8'h5A;
w_real[225] = 8'h5C; w_imag[225] = 8'h58;
w_real[226] = 8'h5E; w_imag[226] = 8'h55;
w_real[227] = 8'h60; w_imag[227] = 8'h53;
w_real[228] = 8'h62; w_imag[228] = 8'h51;
w_real[229] = 8'h64; w_imag[229] = 8'h4E;
w_real[230] = 8'h66; w_imag[230] = 8'h4C;
w_real[231] = 8'h68; w_imag[231] = 8'h49;
w_real[232] = 8'h6A; w_imag[232] = 8'h47;
w_real[233] = 8'h6C; w_imag[233] = 8'h44;
w_real[234] = 8'h6D; w_imag[234] = 8'h41;
w_real[235] = 8'h6F; w_imag[235] = 8'h3F;
w_real[236] = 8'h70; w_imag[236] = 8'h3C;
w_real[237] = 8'h72; w_imag[237] = 8'h39;
w_real[238] = 8'h73; w_imag[238] = 8'h36;
w_real[239] = 8'h75; w_imag[239] = 8'h33;
w_real[240] = 8'h76; w_imag[240] = 8'h30;
w_real[241] = 8'h77; w_imag[241] = 8'h2E;
w_real[242] = 8'h78; w_imag[242] = 8'h2B;
w_real[243] = 8'h79; w_imag[243] = 8'h28;
w_real[244] = 8'h7A; w_imag[244] = 8'h25;
w_real[245] = 8'h7B; w_imag[245] = 8'h22;
w_real[246] = 8'h7C; w_imag[246] = 8'h1F;
w_real[247] = 8'h7C; w_imag[247] = 8'h1C;
w_real[248] = 8'h7D; w_imag[248] = 8'h18;
w_real[249] = 8'h7E; w_imag[249] = 8'h15;
w_real[250] = 8'h7E; w_imag[250] = 8'h12;
w_real[251] = 8'h7F; w_imag[251] = 8'h0F;
w_real[252] = 8'h7F; w_imag[252] = 8'h0C;
w_real[253] = 8'h7F; w_imag[253] = 8'h09;
w_real[254] = 8'h7F; w_imag[254] = 8'h06;
w_real[255] = 8'h7F; w_imag[255] = 8'h03;
