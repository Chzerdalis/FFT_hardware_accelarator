gen_input_real[0] = 16'sd0;
gen_input_real[256] = 16'sd127;
gen_input_real[512] = -16'sd8;
gen_input_real[768] = -16'sd74;
gen_input_real[64] = 16'sd3;
gen_input_real[320] = 16'sd33;
gen_input_real[576] = 16'sd9;
gen_input_real[832] = -16'sd27;
gen_input_real[128] = -16'sd16;
gen_input_real[384] = 16'sd35;
gen_input_real[640] = 16'sd7;
gen_input_real[896] = -16'sd41;
gen_input_real[192] = 16'sd7;
gen_input_real[448] = 16'sd40;
gen_input_real[704] = -16'sd16;
gen_input_real[960] = -16'sd30;
gen_input_real[16] = 16'sd9;
gen_input_real[272] = 16'sd20;
gen_input_real[528] = 16'sd4;
gen_input_real[784] = -16'sd26;
gen_input_real[80] = -16'sd11;
gen_input_real[336] = 16'sd37;
gen_input_real[592] = 16'sd5;
gen_input_real[848] = -16'sd32;
gen_input_real[144] = 16'sd8;
gen_input_real[400] = 16'sd17;
gen_input_real[656] = -16'sd15;
gen_input_real[912] = -16'sd10;
gen_input_real[208] = 16'sd3;
gen_input_real[464] = 16'sd15;
gen_input_real[720] = 16'sd17;
gen_input_real[976] = -16'sd27;
gen_input_real[32] = -16'sd33;
gen_input_real[288] = 16'sd46;
gen_input_real[544] = 16'sd43;
gen_input_real[800] = -16'sd59;
gen_input_real[96] = -16'sd51;
gen_input_real[352] = 16'sd57;
gen_input_real[608] = 16'sd53;
gen_input_real[864] = -16'sd46;
gen_input_real[160] = -16'sd50;
gen_input_real[416] = 16'sd45;
gen_input_real[672] = 16'sd44;
gen_input_real[928] = -16'sd51;
gen_input_real[224] = -16'sd38;
gen_input_real[480] = 16'sd44;
gen_input_real[736] = 16'sd34;
gen_input_real[992] = -16'sd22;
gen_input_real[48] = -16'sd37;
gen_input_real[304] = 16'sd7;
gen_input_real[560] = 16'sd35;
gen_input_real[816] = -16'sd16;
gen_input_real[112] = -16'sd19;
gen_input_real[368] = 16'sd38;
gen_input_real[624] = 16'sd1;
gen_input_real[880] = -16'sd52;
gen_input_real[176] = 16'sd2;
gen_input_real[432] = 16'sd51;
gen_input_real[688] = 16'sd5;
gen_input_real[944] = -16'sd46;
gen_input_real[240] = -16'sd8;
gen_input_real[496] = 16'sd44;
gen_input_real[752] = 16'sd5;
gen_input_real[1008] = -16'sd37;
gen_input_real[4] = -16'sd4;
gen_input_real[260] = 16'sd24;
gen_input_real[516] = 16'sd5;
gen_input_real[772] = -16'sd11;
gen_input_real[68] = -16'sd9;
gen_input_real[324] = 16'sd2;
gen_input_real[580] = 16'sd17;
gen_input_real[836] = -16'sd3;
gen_input_real[132] = -16'sd29;
gen_input_real[388] = 16'sd14;
gen_input_real[644] = 16'sd40;
gen_input_real[900] = -16'sd21;
gen_input_real[196] = -16'sd53;
gen_input_real[452] = 16'sd16;
gen_input_real[708] = 16'sd63;
gen_input_real[964] = -16'sd4;
gen_input_real[20] = -16'sd58;
gen_input_real[276] = -16'sd8;
gen_input_real[532] = 16'sd40;
gen_input_real[788] = 16'sd24;
gen_input_real[84] = -16'sd27;
gen_input_real[340] = -16'sd32;
gen_input_real[596] = 16'sd19;
gen_input_real[852] = 16'sd21;
gen_input_real[148] = -16'sd16;
gen_input_real[404] = 16'sd5;
gen_input_real[660] = 16'sd30;
gen_input_real[916] = -16'sd27;
gen_input_real[212] = -16'sd48;
gen_input_real[468] = 16'sd37;
gen_input_real[724] = 16'sd48;
gen_input_real[980] = -16'sd39;
gen_input_real[36] = -16'sd33;
gen_input_real[292] = 16'sd37;
gen_input_real[548] = 16'sd24;
gen_input_real[804] = -16'sd32;
gen_input_real[100] = -16'sd26;
gen_input_real[356] = 16'sd26;
gen_input_real[612] = 16'sd29;
gen_input_real[868] = -16'sd26;
gen_input_real[164] = -16'sd26;
gen_input_real[420] = 16'sd29;
gen_input_real[676] = 16'sd13;
gen_input_real[932] = -16'sd20;
gen_input_real[228] = -16'sd3;
gen_input_real[484] = 16'sd2;
gen_input_real[740] = 16'sd14;
gen_input_real[996] = 16'sd8;
gen_input_real[52] = -16'sd39;
gen_input_real[308] = -16'sd10;
gen_input_real[564] = 16'sd43;
gen_input_real[820] = 16'sd6;
gen_input_real[116] = -16'sd18;
gen_input_real[372] = -16'sd4;
gen_input_real[628] = -16'sd8;
gen_input_real[884] = 16'sd9;
gen_input_real[180] = 16'sd16;
gen_input_real[436] = -16'sd23;
gen_input_real[692] = -16'sd10;
gen_input_real[948] = 16'sd34;
gen_input_real[244] = 16'sd3;
gen_input_real[500] = -16'sd33;
gen_input_real[756] = 16'sd4;
gen_input_real[1012] = 16'sd23;
gen_input_real[8] = -16'sd10;
gen_input_real[264] = -16'sd11;
gen_input_real[520] = 16'sd14;
gen_input_real[776] = 16'sd0;
gen_input_real[72] = -16'sd21;
gen_input_real[328] = 16'sd12;
gen_input_real[584] = 16'sd36;
gen_input_real[840] = -16'sd17;
gen_input_real[136] = -16'sd51;
gen_input_real[392] = 16'sd10;
gen_input_real[648] = 16'sd54;
gen_input_real[904] = 16'sd1;
gen_input_real[200] = -16'sd45;
gen_input_real[456] = -16'sd9;
gen_input_real[712] = 16'sd28;
gen_input_real[968] = 16'sd9;
gen_input_real[24] = -16'sd14;
gen_input_real[280] = -16'sd6;
gen_input_real[536] = 16'sd10;
gen_input_real[792] = 16'sd1;
gen_input_real[88] = -16'sd15;
gen_input_real[344] = 16'sd1;
gen_input_real[600] = 16'sd17;
gen_input_real[856] = -16'sd2;
gen_input_real[152] = -16'sd16;
gen_input_real[408] = 16'sd7;
gen_input_real[664] = 16'sd12;
gen_input_real[920] = -16'sd14;
gen_input_real[216] = -16'sd4;
gen_input_real[472] = 16'sd17;
gen_input_real[728] = -16'sd13;
gen_input_real[984] = -16'sd9;
gen_input_real[40] = 16'sd44;
gen_input_real[296] = -16'sd2;
gen_input_real[552] = -16'sd62;
gen_input_real[808] = 16'sd6;
gen_input_real[104] = 16'sd42;
gen_input_real[360] = 16'sd6;
gen_input_real[616] = -16'sd7;
gen_input_real[872] = -16'sd23;
gen_input_real[168] = -16'sd10;
gen_input_real[424] = 16'sd20;
gen_input_real[680] = 16'sd12;
gen_input_real[936] = 16'sd0;
gen_input_real[232] = -16'sd13;
gen_input_real[488] = -16'sd18;
gen_input_real[744] = 16'sd15;
gen_input_real[1000] = 16'sd27;
gen_input_real[56] = -16'sd12;
gen_input_real[312] = -16'sd25;
gen_input_real[568] = 16'sd7;
gen_input_real[824] = 16'sd14;
gen_input_real[120] = -16'sd1;
gen_input_real[376] = -16'sd8;
gen_input_real[632] = -16'sd7;
gen_input_real[888] = 16'sd17;
gen_input_real[184] = 16'sd7;
gen_input_real[440] = -16'sd26;
gen_input_real[696] = 16'sd5;
gen_input_real[952] = 16'sd20;
gen_input_real[248] = -16'sd14;
gen_input_real[504] = -16'sd3;
gen_input_real[760] = 16'sd16;
gen_input_real[1016] = -16'sd13;
gen_input_real[12] = -16'sd14;
gen_input_real[268] = 16'sd27;
gen_input_real[524] = 16'sd7;
gen_input_real[780] = -16'sd35;
gen_input_real[76] = 16'sd5;
gen_input_real[332] = 16'sd36;
gen_input_real[588] = -16'sd14;
gen_input_real[844] = -16'sd39;
gen_input_real[140] = 16'sd9;
gen_input_real[396] = 16'sd44;
gen_input_real[652] = 16'sd0;
gen_input_real[908] = -16'sd41;
gen_input_real[204] = 16'sd2;
gen_input_real[460] = 16'sd27;
gen_input_real[716] = -16'sd7;
gen_input_real[972] = -16'sd16;
gen_input_real[28] = 16'sd0;
gen_input_real[284] = 16'sd21;
gen_input_real[540] = 16'sd14;
gen_input_real[796] = -16'sd32;
gen_input_real[92] = -16'sd15;
gen_input_real[348] = 16'sd25;
gen_input_real[604] = -16'sd2;
gen_input_real[860] = -16'sd2;
gen_input_real[156] = 16'sd23;
gen_input_real[412] = -16'sd14;
gen_input_real[668] = -16'sd36;
gen_input_real[924] = 16'sd12;
gen_input_real[220] = 16'sd40;
gen_input_real[476] = 16'sd0;
gen_input_real[732] = -16'sd36;
gen_input_real[988] = -16'sd12;
gen_input_real[44] = 16'sd26;
gen_input_real[300] = 16'sd19;
gen_input_real[556] = -16'sd13;
gen_input_real[812] = -16'sd16;
gen_input_real[108] = -16'sd2;
gen_input_real[364] = 16'sd7;
gen_input_real[620] = 16'sd19;
gen_input_real[876] = -16'sd6;
gen_input_real[172] = -16'sd31;
gen_input_real[428] = 16'sd17;
gen_input_real[684] = 16'sd29;
gen_input_real[940] = -16'sd32;
gen_input_real[236] = -16'sd16;
gen_input_real[492] = 16'sd40;
gen_input_real[748] = 16'sd5;
gen_input_real[1004] = -16'sd40;
gen_input_real[60] = -16'sd5;
gen_input_real[316] = 16'sd32;
gen_input_real[572] = 16'sd18;
gen_input_real[828] = -16'sd19;
gen_input_real[124] = -16'sd40;
gen_input_real[380] = 16'sd19;
gen_input_real[636] = 16'sd61;
gen_input_real[892] = -16'sd33;
gen_input_real[188] = -16'sd56;
gen_input_real[444] = 16'sd34;
gen_input_real[700] = 16'sd20;
gen_input_real[956] = -16'sd19;
gen_input_real[252] = 16'sd12;
gen_input_real[508] = 16'sd19;
gen_input_real[764] = -16'sd20;
gen_input_real[1020] = -16'sd40;
gen_input_real[1] = 16'sd12;
gen_input_real[257] = 16'sd56;
gen_input_real[513] = -16'sd6;
gen_input_real[769] = -16'sd58;
gen_input_real[65] = 16'sd9;
gen_input_real[321] = 16'sd55;
gen_input_real[577] = -16'sd16;
gen_input_real[833] = -16'sd44;
gen_input_real[129] = 16'sd14;
gen_input_real[385] = 16'sd26;
gen_input_real[641] = 16'sd0;
gen_input_real[897] = -16'sd19;
gen_input_real[193] = -16'sd23;
gen_input_real[449] = 16'sd24;
gen_input_real[705] = 16'sd40;
gen_input_real[961] = -16'sd30;
gen_input_real[17] = -16'sd35;
gen_input_real[273] = 16'sd33;
gen_input_real[529] = 16'sd17;
gen_input_real[785] = -16'sd29;
gen_input_real[81] = -16'sd10;
gen_input_real[337] = 16'sd10;
gen_input_real[593] = 16'sd19;
gen_input_real[849] = 16'sd9;
gen_input_real[145] = -16'sd32;
gen_input_real[401] = -16'sd10;
gen_input_real[657] = 16'sd40;
gen_input_real[913] = -16'sd2;
gen_input_real[209] = -16'sd44;
gen_input_real[465] = 16'sd7;
gen_input_real[721] = 16'sd42;
gen_input_real[977] = -16'sd5;
gen_input_real[33] = -16'sd38;
gen_input_real[289] = 16'sd9;
gen_input_real[545] = 16'sd43;
gen_input_real[801] = -16'sd23;
gen_input_real[97] = -16'sd47;
gen_input_real[353] = 16'sd35;
gen_input_real[609] = 16'sd35;
gen_input_real[865] = -16'sd43;
gen_input_real[161] = -16'sd18;
gen_input_real[417] = 16'sd52;
gen_input_real[673] = 16'sd16;
gen_input_real[929] = -16'sd61;
gen_input_real[225] = -16'sd30;
gen_input_real[481] = 16'sd63;
gen_input_real[737] = 16'sd49;
gen_input_real[993] = -16'sd51;
gen_input_real[49] = -16'sd63;
gen_input_real[305] = 16'sd29;
gen_input_real[561] = 16'sd66;
gen_input_real[817] = -16'sd11;
gen_input_real[113] = -16'sd54;
gen_input_real[369] = 16'sd11;
gen_input_real[625] = 16'sd36;
gen_input_real[881] = -16'sd21;
gen_input_real[177] = -16'sd24;
gen_input_real[433] = 16'sd23;
gen_input_real[689] = 16'sd19;
gen_input_real[945] = -16'sd18;
gen_input_real[241] = -16'sd13;
gen_input_real[497] = 16'sd13;
gen_input_real[753] = 16'sd9;
gen_input_real[1009] = -16'sd4;
gen_input_real[5] = -16'sd15;
gen_input_real[261] = -16'sd10;
gen_input_real[517] = 16'sd28;
gen_input_real[773] = 16'sd23;
gen_input_real[69] = -16'sd38;
gen_input_real[325] = -16'sd26;
gen_input_real[581] = 16'sd40;
gen_input_real[837] = 16'sd15;
gen_input_real[133] = -16'sd32;
gen_input_real[389] = 16'sd2;
gen_input_real[645] = 16'sd27;
gen_input_real[901] = -16'sd15;
gen_input_real[197] = -16'sd36;
gen_input_real[453] = 16'sd20;
gen_input_real[709] = 16'sd54;
gen_input_real[965] = -16'sd20;
gen_input_real[21] = -16'sd66;
gen_input_real[277] = 16'sd13;
gen_input_real[533] = 16'sd77;
gen_input_real[789] = 16'sd1;
gen_input_real[85] = -16'sd81;
gen_input_real[341] = -16'sd13;
gen_input_real[597] = 16'sd73;
gen_input_real[853] = 16'sd16;
gen_input_real[149] = -16'sd62;
gen_input_real[405] = -16'sd12;
gen_input_real[661] = 16'sd64;
gen_input_real[917] = 16'sd7;
gen_input_real[213] = -16'sd68;
gen_input_real[469] = -16'sd6;
gen_input_real[725] = 16'sd61;
gen_input_real[981] = 16'sd0;
gen_input_real[37] = -16'sd47;
gen_input_real[293] = 16'sd13;
gen_input_real[549] = 16'sd27;
gen_input_real[805] = -16'sd23;
gen_input_real[101] = -16'sd4;
gen_input_real[357] = 16'sd15;
gen_input_real[613] = 16'sd0;
gen_input_real[869] = 16'sd4;
gen_input_real[165] = -16'sd21;
gen_input_real[421] = -16'sd16;
gen_input_real[677] = 16'sd37;
gen_input_real[933] = 16'sd9;
gen_input_real[229] = -16'sd33;
gen_input_real[485] = 16'sd2;
gen_input_real[741] = 16'sd27;
gen_input_real[997] = -16'sd4;
gen_input_real[53] = -16'sd30;
gen_input_real[309] = -16'sd9;
gen_input_real[565] = 16'sd30;
gen_input_real[821] = 16'sd22;
gen_input_real[117] = -16'sd26;
gen_input_real[373] = -16'sd22;
gen_input_real[629] = 16'sd34;
gen_input_real[885] = 16'sd19;
gen_input_real[181] = -16'sd47;
gen_input_real[437] = -16'sd25;
gen_input_real[693] = 16'sd48;
gen_input_real[949] = 16'sd40;
gen_input_real[245] = -16'sd45;
gen_input_real[501] = -16'sd61;
gen_input_real[757] = 16'sd47;
gen_input_real[1013] = 16'sd80;
gen_input_real[9] = -16'sd48;
gen_input_real[265] = -16'sd76;
gen_input_real[521] = 16'sd39;
gen_input_real[777] = 16'sd49;
gen_input_real[73] = -16'sd31;
gen_input_real[329] = -16'sd17;
gen_input_real[585] = 16'sd28;
gen_input_real[841] = -16'sd3;
gen_input_real[137] = -16'sd28;
gen_input_real[393] = 16'sd8;
gen_input_real[649] = 16'sd33;
gen_input_real[905] = -16'sd1;
gen_input_real[201] = -16'sd41;
gen_input_real[457] = -16'sd12;
gen_input_real[713] = 16'sd41;
gen_input_real[969] = 16'sd21;
gen_input_real[25] = -16'sd32;
gen_input_real[281] = -16'sd19;
gen_input_real[537] = 16'sd31;
gen_input_real[793] = 16'sd16;
gen_input_real[89] = -16'sd40;
gen_input_real[345] = -16'sd12;
gen_input_real[601] = 16'sd40;
gen_input_real[857] = 16'sd0;
gen_input_real[153] = -16'sd22;
gen_input_real[409] = 16'sd6;
gen_input_real[665] = 16'sd9;
gen_input_real[921] = 16'sd7;
gen_input_real[217] = -16'sd16;
gen_input_real[473] = -16'sd32;
gen_input_real[729] = 16'sd26;
gen_input_real[985] = 16'sd44;
gen_input_real[41] = -16'sd15;
gen_input_real[297] = -16'sd47;
gen_input_real[553] = -16'sd13;
gen_input_real[809] = 16'sd53;
gen_input_real[105] = 16'sd31;
gen_input_real[361] = -16'sd55;
gen_input_real[617] = -16'sd26;
gen_input_real[873] = 16'sd53;
gen_input_real[169] = 16'sd8;
gen_input_real[425] = -16'sd49;
gen_input_real[681] = 16'sd12;
gen_input_real[937] = 16'sd37;
gen_input_real[233] = -16'sd20;
gen_input_real[489] = -16'sd15;
gen_input_real[745] = 16'sd10;
gen_input_real[1001] = 16'sd7;
gen_input_real[57] = 16'sd1;
gen_input_real[313] = -16'sd20;
gen_input_real[569] = 16'sd4;
gen_input_real[825] = 16'sd34;
gen_input_real[121] = -16'sd24;
gen_input_real[377] = -16'sd39;
gen_input_real[633] = 16'sd42;
gen_input_real[889] = 16'sd40;
gen_input_real[185] = -16'sd47;
gen_input_real[441] = -16'sd37;
gen_input_real[697] = 16'sd38;
gen_input_real[953] = 16'sd34;
gen_input_real[249] = -16'sd23;
gen_input_real[505] = -16'sd33;
gen_input_real[761] = 16'sd16;
gen_input_real[1017] = 16'sd27;
gen_input_real[13] = -16'sd23;
gen_input_real[269] = -16'sd12;
gen_input_real[525] = 16'sd24;
gen_input_real[781] = -16'sd1;
gen_input_real[77] = -16'sd5;
gen_input_real[333] = 16'sd0;
gen_input_real[589] = -16'sd20;
gen_input_real[845] = 16'sd12;
gen_input_real[141] = 16'sd26;
gen_input_real[397] = -16'sd24;
gen_input_real[653] = -16'sd12;
gen_input_real[909] = 16'sd25;
gen_input_real[205] = 16'sd10;
gen_input_real[461] = -16'sd15;
gen_input_real[717] = -16'sd29;
gen_input_real[973] = 16'sd2;
gen_input_real[29] = 16'sd42;
gen_input_real[285] = 16'sd6;
gen_input_real[541] = -16'sd28;
gen_input_real[797] = -16'sd10;
gen_input_real[93] = 16'sd0;
gen_input_real[349] = 16'sd10;
gen_input_real[605] = 16'sd17;
gen_input_real[861] = -16'sd1;
gen_input_real[157] = -16'sd14;
gen_input_real[413] = -16'sd18;
gen_input_real[669] = -16'sd4;
gen_input_real[925] = 16'sd42;
gen_input_real[221] = 16'sd22;
gen_input_real[477] = -16'sd60;
gen_input_real[733] = -16'sd19;
gen_input_real[989] = 16'sd64;
gen_input_real[45] = 16'sd1;
gen_input_real[301] = -16'sd52;
gen_input_real[557] = 16'sd12;
gen_input_real[813] = 16'sd29;
gen_input_real[109] = -16'sd11;
gen_input_real[365] = -16'sd9;
gen_input_real[621] = 16'sd6;
gen_input_real[877] = 16'sd8;
gen_input_real[173] = -16'sd2;
gen_input_real[429] = -16'sd18;
gen_input_real[685] = 16'sd0;
gen_input_real[941] = 16'sd21;
gen_input_real[237] = -16'sd2;
gen_input_real[493] = -16'sd10;
gen_input_real[749] = 16'sd6;
gen_input_real[1005] = -16'sd5;
gen_input_real[61] = 16'sd0;
gen_input_real[317] = 16'sd16;
gen_input_real[573] = -16'sd14;
gen_input_real[829] = -16'sd18;
gen_input_real[125] = 16'sd10;
gen_input_real[381] = 16'sd17;
gen_input_real[637] = 16'sd16;
gen_input_real[893] = -16'sd20;
gen_input_real[189] = -16'sd37;
gen_input_real[445] = 16'sd21;
gen_input_real[701] = 16'sd33;
gen_input_real[957] = -16'sd20;
gen_input_real[253] = -16'sd14;
gen_input_real[509] = 16'sd19;
gen_input_real[765] = -16'sd3;
gen_input_real[1021] = -16'sd16;
gen_input_real[2] = 16'sd16;
gen_input_real[258] = 16'sd3;
gen_input_real[514] = -16'sd19;
gen_input_real[770] = 16'sd14;
gen_input_real[66] = 16'sd20;
gen_input_real[322] = -16'sd33;
gen_input_real[578] = -16'sd21;
gen_input_real[834] = 16'sd37;
gen_input_real[130] = 16'sd20;
gen_input_real[386] = -16'sd16;
gen_input_real[642] = -16'sd17;
gen_input_real[898] = -16'sd10;
gen_input_real[194] = 16'sd18;
gen_input_real[450] = 16'sd14;
gen_input_real[706] = -16'sd16;
gen_input_real[962] = 16'sd0;
gen_input_real[18] = 16'sd5;
gen_input_real[274] = -16'sd6;
gen_input_real[530] = 16'sd10;
gen_input_real[786] = 16'sd2;
gen_input_real[82] = -16'sd21;
gen_input_real[338] = 16'sd0;
gen_input_real[594] = 16'sd18;
gen_input_real[850] = 16'sd2;
gen_input_real[146] = -16'sd8;
gen_input_real[402] = -16'sd6;
gen_input_real[658] = 16'sd9;
gen_input_real[914] = 16'sd11;
gen_input_real[210] = -16'sd29;
gen_input_real[466] = -16'sd12;
gen_input_real[722] = 16'sd52;
gen_input_real[978] = -16'sd1;
gen_input_real[34] = -16'sd64;
gen_input_real[290] = 16'sd19;
gen_input_real[546] = 16'sd60;
gen_input_real[802] = -16'sd22;
gen_input_real[98] = -16'sd42;
gen_input_real[354] = 16'sd4;
gen_input_real[610] = 16'sd18;
gen_input_real[866] = 16'sd14;
gen_input_real[162] = 16'sd1;
gen_input_real[418] = -16'sd17;
gen_input_real[674] = -16'sd10;
gen_input_real[930] = 16'sd0;
gen_input_real[226] = 16'sd10;
gen_input_real[482] = 16'sd28;
gen_input_real[738] = -16'sd6;
gen_input_real[994] = -16'sd42;
gen_input_real[50] = -16'sd2;
gen_input_real[306] = 16'sd29;
gen_input_real[562] = 16'sd15;
gen_input_real[818] = -16'sd10;
gen_input_real[114] = -16'sd25;
gen_input_real[370] = 16'sd12;
gen_input_real[626] = 16'sd24;
gen_input_real[882] = -16'sd26;
gen_input_real[178] = -16'sd12;
gen_input_real[434] = 16'sd20;
gen_input_real[690] = 16'sd0;
gen_input_real[946] = 16'sd5;
gen_input_real[242] = 16'sd1;
gen_input_real[498] = -16'sd24;
gen_input_real[754] = 16'sd12;
gen_input_real[1010] = 16'sd23;
gen_input_real[6] = -16'sd27;
gen_input_real[262] = -16'sd16;
gen_input_real[518] = 16'sd33;
gen_input_real[774] = 16'sd23;
gen_input_real[70] = -16'sd34;
gen_input_real[326] = -16'sd38;
gen_input_real[582] = 16'sd37;
gen_input_real[838] = 16'sd47;
gen_input_real[134] = -16'sd40;
gen_input_real[390] = -16'sd42;
gen_input_real[646] = 16'sd39;
gen_input_real[902] = 16'sd24;
gen_input_real[198] = -16'sd34;
gen_input_real[454] = -16'sd4;
gen_input_real[710] = 16'sd20;
gen_input_real[966] = -16'sd1;
gen_input_real[22] = -16'sd7;
gen_input_real[278] = -16'sd10;
gen_input_real[534] = 16'sd15;
gen_input_real[790] = 16'sd20;
gen_input_real[86] = -16'sd37;
gen_input_real[342] = -16'sd12;
gen_input_real[598] = 16'sd49;
gen_input_real[854] = -16'sd8;
gen_input_real[150] = -16'sd53;
gen_input_real[406] = 16'sd26;
gen_input_real[662] = 16'sd55;
gen_input_real[918] = -16'sd31;
gen_input_real[214] = -16'sd53;
gen_input_real[470] = 16'sd13;
gen_input_real[726] = 16'sd47;
gen_input_real[982] = 16'sd15;
gen_input_real[38] = -16'sd44;
gen_input_real[294] = -16'sd26;
gen_input_real[550] = 16'sd32;
gen_input_real[806] = 16'sd16;
gen_input_real[102] = -16'sd7;
gen_input_real[358] = -16'sd9;
gen_input_real[614] = -16'sd6;
gen_input_real[870] = 16'sd22;
gen_input_real[166] = 16'sd0;
gen_input_real[422] = -16'sd40;
gen_input_real[678] = 16'sd12;
gen_input_real[934] = 16'sd40;
gen_input_real[230] = -16'sd16;
gen_input_real[486] = -16'sd31;
gen_input_real[742] = 16'sd19;
gen_input_real[998] = 16'sd32;
gen_input_real[54] = -16'sd21;
gen_input_real[310] = -16'sd41;
gen_input_real[566] = 16'sd12;
gen_input_real[822] = 16'sd41;
gen_input_real[118] = 16'sd1;
gen_input_real[374] = -16'sd33;
gen_input_real[630] = -16'sd8;
gen_input_real[886] = 16'sd28;
gen_input_real[182] = 16'sd3;
gen_input_real[438] = -16'sd28;
gen_input_real[694] = 16'sd17;
gen_input_real[950] = 16'sd31;
gen_input_real[246] = -16'sd49;
gen_input_real[502] = -16'sd39;
gen_input_real[758] = 16'sd76;
gen_input_real[1014] = 16'sd48;
gen_input_real[10] = -16'sd80;
gen_input_real[266] = -16'sd47;
gen_input_real[522] = 16'sd61;
gen_input_real[778] = 16'sd45;
gen_input_real[74] = -16'sd40;
gen_input_real[330] = -16'sd48;
gen_input_real[586] = 16'sd25;
gen_input_real[842] = 16'sd47;
gen_input_real[138] = -16'sd19;
gen_input_real[394] = -16'sd34;
gen_input_real[650] = 16'sd22;
gen_input_real[906] = 16'sd26;
gen_input_real[202] = -16'sd22;
gen_input_real[458] = -16'sd30;
gen_input_real[714] = 16'sd9;
gen_input_real[970] = 16'sd30;
gen_input_real[26] = 16'sd4;
gen_input_real[282] = -16'sd27;
gen_input_real[538] = -16'sd2;
gen_input_real[794] = 16'sd33;
gen_input_real[90] = -16'sd9;
gen_input_real[346] = -16'sd37;
gen_input_real[602] = 16'sd16;
gen_input_real[858] = 16'sd21;
gen_input_real[154] = -16'sd4;
gen_input_real[410] = 16'sd0;
gen_input_real[666] = -16'sd15;
gen_input_real[922] = 16'sd4;
gen_input_real[218] = 16'sd23;
gen_input_real[474] = -16'sd27;
gen_input_real[730] = -16'sd13;
gen_input_real[986] = 16'sd47;
gen_input_real[42] = 16'sd0;
gen_input_real[298] = -16'sd61;
gen_input_real[554] = 16'sd6;
gen_input_real[810] = 16'sd68;
gen_input_real[106] = -16'sd7;
gen_input_real[362] = -16'sd64;
gen_input_real[618] = 16'sd12;
gen_input_real[874] = 16'sd62;
gen_input_real[170] = -16'sd16;
gen_input_real[426] = -16'sd73;
gen_input_real[682] = 16'sd13;
gen_input_real[938] = 16'sd81;
gen_input_real[234] = -16'sd1;
gen_input_real[490] = -16'sd77;
gen_input_real[746] = -16'sd13;
gen_input_real[1002] = 16'sd66;
gen_input_real[58] = 16'sd20;
gen_input_real[314] = -16'sd54;
gen_input_real[570] = -16'sd20;
gen_input_real[826] = 16'sd36;
gen_input_real[122] = 16'sd15;
gen_input_real[378] = -16'sd27;
gen_input_real[634] = -16'sd2;
gen_input_real[890] = 16'sd32;
gen_input_real[186] = -16'sd15;
gen_input_real[442] = -16'sd40;
gen_input_real[698] = 16'sd26;
gen_input_real[954] = 16'sd38;
gen_input_real[250] = -16'sd23;
gen_input_real[506] = -16'sd28;
gen_input_real[762] = 16'sd10;
gen_input_real[1018] = 16'sd15;
gen_input_real[14] = 16'sd4;
gen_input_real[270] = -16'sd9;
gen_input_real[526] = -16'sd13;
gen_input_real[782] = 16'sd13;
gen_input_real[78] = 16'sd18;
gen_input_real[334] = -16'sd19;
gen_input_real[590] = -16'sd23;
gen_input_real[846] = 16'sd24;
gen_input_real[142] = 16'sd21;
gen_input_real[398] = -16'sd36;
gen_input_real[654] = -16'sd11;
gen_input_real[910] = 16'sd54;
gen_input_real[206] = 16'sd11;
gen_input_real[462] = -16'sd66;
gen_input_real[718] = -16'sd29;
gen_input_real[974] = 16'sd63;
gen_input_real[30] = 16'sd51;
gen_input_real[286] = -16'sd49;
gen_input_real[542] = -16'sd63;
gen_input_real[798] = 16'sd30;
gen_input_real[94] = 16'sd61;
gen_input_real[350] = -16'sd16;
gen_input_real[606] = -16'sd52;
gen_input_real[862] = 16'sd18;
gen_input_real[158] = 16'sd43;
gen_input_real[414] = -16'sd35;
gen_input_real[670] = -16'sd35;
gen_input_real[926] = 16'sd47;
gen_input_real[222] = 16'sd23;
gen_input_real[478] = -16'sd43;
gen_input_real[734] = -16'sd9;
gen_input_real[990] = 16'sd38;
gen_input_real[46] = 16'sd5;
gen_input_real[302] = -16'sd42;
gen_input_real[558] = -16'sd7;
gen_input_real[814] = 16'sd44;
gen_input_real[110] = 16'sd2;
gen_input_real[366] = -16'sd40;
gen_input_real[622] = 16'sd10;
gen_input_real[878] = 16'sd32;
gen_input_real[174] = -16'sd9;
gen_input_real[430] = -16'sd19;
gen_input_real[686] = -16'sd10;
gen_input_real[942] = 16'sd10;
gen_input_real[238] = 16'sd29;
gen_input_real[494] = -16'sd17;
gen_input_real[750] = -16'sd33;
gen_input_real[1006] = 16'sd35;
gen_input_real[62] = 16'sd30;
gen_input_real[318] = -16'sd40;
gen_input_real[574] = -16'sd24;
gen_input_real[830] = 16'sd23;
gen_input_real[126] = 16'sd19;
gen_input_real[382] = 16'sd0;
gen_input_real[638] = -16'sd26;
gen_input_real[894] = -16'sd14;
gen_input_real[190] = 16'sd44;
gen_input_real[446] = 16'sd16;
gen_input_real[702] = -16'sd55;
gen_input_real[958] = -16'sd9;
gen_input_real[254] = 16'sd58;
gen_input_real[510] = 16'sd6;
gen_input_real[766] = -16'sd56;
gen_input_real[1022] = -16'sd12;
gen_input_real[3] = 16'sd40;
gen_input_real[259] = 16'sd20;
gen_input_real[515] = -16'sd19;
gen_input_real[771] = -16'sd12;
gen_input_real[67] = 16'sd19;
gen_input_real[323] = -16'sd20;
gen_input_real[579] = -16'sd34;
gen_input_real[835] = 16'sd56;
gen_input_real[131] = 16'sd33;
gen_input_real[387] = -16'sd61;
gen_input_real[643] = -16'sd19;
gen_input_real[899] = 16'sd40;
gen_input_real[195] = 16'sd19;
gen_input_real[451] = -16'sd18;
gen_input_real[707] = -16'sd32;
gen_input_real[963] = 16'sd5;
gen_input_real[19] = 16'sd40;
gen_input_real[275] = -16'sd5;
gen_input_real[531] = -16'sd40;
gen_input_real[787] = 16'sd16;
gen_input_real[83] = 16'sd32;
gen_input_real[339] = -16'sd29;
gen_input_real[595] = -16'sd17;
gen_input_real[851] = 16'sd31;
gen_input_real[147] = 16'sd6;
gen_input_real[403] = -16'sd19;
gen_input_real[659] = -16'sd7;
gen_input_real[915] = 16'sd2;
gen_input_real[211] = 16'sd16;
gen_input_real[467] = 16'sd13;
gen_input_real[723] = -16'sd19;
gen_input_real[979] = -16'sd26;
gen_input_real[35] = 16'sd12;
gen_input_real[291] = 16'sd36;
gen_input_real[547] = 16'sd0;
gen_input_real[803] = -16'sd40;
gen_input_real[99] = -16'sd12;
gen_input_real[355] = 16'sd36;
gen_input_real[611] = 16'sd14;
gen_input_real[867] = -16'sd23;
gen_input_real[163] = 16'sd2;
gen_input_real[419] = 16'sd2;
gen_input_real[675] = -16'sd25;
gen_input_real[931] = 16'sd15;
gen_input_real[227] = 16'sd32;
gen_input_real[483] = -16'sd14;
gen_input_real[739] = -16'sd21;
gen_input_real[995] = 16'sd0;
gen_input_real[51] = 16'sd16;
gen_input_real[307] = 16'sd7;
gen_input_real[563] = -16'sd27;
gen_input_real[819] = -16'sd2;
gen_input_real[115] = 16'sd41;
gen_input_real[371] = 16'sd0;
gen_input_real[627] = -16'sd44;
gen_input_real[883] = -16'sd9;
gen_input_real[179] = 16'sd39;
gen_input_real[435] = 16'sd14;
gen_input_real[691] = -16'sd36;
gen_input_real[947] = -16'sd5;
gen_input_real[243] = 16'sd35;
gen_input_real[499] = -16'sd7;
gen_input_real[755] = -16'sd27;
gen_input_real[1011] = 16'sd14;
gen_input_real[7] = 16'sd13;
gen_input_real[263] = -16'sd16;
gen_input_real[519] = 16'sd3;
gen_input_real[775] = 16'sd14;
gen_input_real[71] = -16'sd20;
gen_input_real[327] = -16'sd5;
gen_input_real[583] = 16'sd26;
gen_input_real[839] = -16'sd7;
gen_input_real[135] = -16'sd17;
gen_input_real[391] = 16'sd7;
gen_input_real[647] = 16'sd8;
gen_input_real[903] = 16'sd1;
gen_input_real[199] = -16'sd14;
gen_input_real[455] = -16'sd7;
gen_input_real[711] = 16'sd25;
gen_input_real[967] = 16'sd12;
gen_input_real[23] = -16'sd27;
gen_input_real[279] = -16'sd15;
gen_input_real[535] = 16'sd18;
gen_input_real[791] = 16'sd13;
gen_input_real[87] = 16'sd0;
gen_input_real[343] = -16'sd12;
gen_input_real[599] = -16'sd20;
gen_input_real[855] = 16'sd10;
gen_input_real[151] = 16'sd23;
gen_input_real[407] = 16'sd7;
gen_input_real[663] = -16'sd6;
gen_input_real[919] = -16'sd42;
gen_input_real[215] = -16'sd6;
gen_input_real[471] = 16'sd62;
gen_input_real[727] = 16'sd2;
gen_input_real[983] = -16'sd44;
gen_input_real[39] = 16'sd9;
gen_input_real[295] = 16'sd13;
gen_input_real[551] = -16'sd17;
gen_input_real[807] = 16'sd4;
gen_input_real[103] = 16'sd14;
gen_input_real[359] = -16'sd12;
gen_input_real[615] = -16'sd7;
gen_input_real[871] = 16'sd16;
gen_input_real[167] = 16'sd2;
gen_input_real[423] = -16'sd17;
gen_input_real[679] = -16'sd1;
gen_input_real[935] = 16'sd15;
gen_input_real[231] = -16'sd1;
gen_input_real[487] = -16'sd10;
gen_input_real[743] = 16'sd6;
gen_input_real[999] = 16'sd14;
gen_input_real[55] = -16'sd9;
gen_input_real[311] = -16'sd28;
gen_input_real[567] = 16'sd9;
gen_input_real[823] = 16'sd45;
gen_input_real[119] = -16'sd1;
gen_input_real[375] = -16'sd54;
gen_input_real[631] = -16'sd10;
gen_input_real[887] = 16'sd51;
gen_input_real[183] = 16'sd17;
gen_input_real[439] = -16'sd36;
gen_input_real[695] = -16'sd12;
gen_input_real[951] = 16'sd21;
gen_input_real[247] = 16'sd0;
gen_input_real[503] = -16'sd14;
gen_input_real[759] = 16'sd11;
gen_input_real[1015] = 16'sd10;
gen_input_real[11] = -16'sd23;
gen_input_real[267] = -16'sd4;
gen_input_real[523] = 16'sd33;
gen_input_real[779] = -16'sd3;
gen_input_real[75] = -16'sd34;
gen_input_real[331] = 16'sd10;
gen_input_real[587] = 16'sd23;
gen_input_real[843] = -16'sd16;
gen_input_real[139] = -16'sd9;
gen_input_real[395] = 16'sd8;
gen_input_real[651] = 16'sd4;
gen_input_real[907] = 16'sd18;
gen_input_real[203] = -16'sd6;
gen_input_real[459] = -16'sd43;
gen_input_real[715] = 16'sd10;
gen_input_real[971] = 16'sd39;
gen_input_real[27] = -16'sd8;
gen_input_real[283] = -16'sd14;
gen_input_real[539] = -16'sd2;
gen_input_real[795] = 16'sd3;
gen_input_real[91] = 16'sd20;
gen_input_real[347] = -16'sd13;
gen_input_real[603] = -16'sd29;
gen_input_real[859] = 16'sd26;
gen_input_real[155] = 16'sd26;
gen_input_real[411] = -16'sd29;
gen_input_real[667] = -16'sd26;
gen_input_real[923] = 16'sd26;
gen_input_real[219] = 16'sd32;
gen_input_real[475] = -16'sd24;
gen_input_real[731] = -16'sd37;
gen_input_real[987] = 16'sd33;
gen_input_real[43] = 16'sd39;
gen_input_real[299] = -16'sd48;
gen_input_real[555] = -16'sd37;
gen_input_real[811] = 16'sd48;
gen_input_real[107] = 16'sd27;
gen_input_real[363] = -16'sd30;
gen_input_real[619] = -16'sd5;
gen_input_real[875] = 16'sd16;
gen_input_real[171] = -16'sd21;
gen_input_real[427] = -16'sd19;
gen_input_real[683] = 16'sd32;
gen_input_real[939] = 16'sd27;
gen_input_real[235] = -16'sd24;
gen_input_real[491] = -16'sd40;
gen_input_real[747] = 16'sd8;
gen_input_real[1003] = 16'sd58;
gen_input_real[59] = 16'sd4;
gen_input_real[315] = -16'sd63;
gen_input_real[571] = -16'sd16;
gen_input_real[827] = 16'sd53;
gen_input_real[123] = 16'sd21;
gen_input_real[379] = -16'sd40;
gen_input_real[635] = -16'sd14;
gen_input_real[891] = 16'sd29;
gen_input_real[187] = 16'sd3;
gen_input_real[443] = -16'sd17;
gen_input_real[699] = -16'sd2;
gen_input_real[955] = 16'sd9;
gen_input_real[251] = 16'sd11;
gen_input_real[507] = -16'sd5;
gen_input_real[763] = -16'sd24;
gen_input_real[1019] = 16'sd4;
gen_input_real[15] = 16'sd37;
gen_input_real[271] = -16'sd5;
gen_input_real[527] = -16'sd44;
gen_input_real[783] = 16'sd8;
gen_input_real[79] = 16'sd46;
gen_input_real[335] = -16'sd5;
gen_input_real[591] = -16'sd51;
gen_input_real[847] = -16'sd2;
gen_input_real[143] = 16'sd52;
gen_input_real[399] = -16'sd1;
gen_input_real[655] = -16'sd38;
gen_input_real[911] = 16'sd19;
gen_input_real[207] = 16'sd16;
gen_input_real[463] = -16'sd35;
gen_input_real[719] = -16'sd7;
gen_input_real[975] = 16'sd37;
gen_input_real[31] = 16'sd22;
gen_input_real[287] = -16'sd34;
gen_input_real[543] = -16'sd44;
gen_input_real[799] = 16'sd38;
gen_input_real[95] = 16'sd51;
gen_input_real[351] = -16'sd44;
gen_input_real[607] = -16'sd45;
gen_input_real[863] = 16'sd50;
gen_input_real[159] = 16'sd46;
gen_input_real[415] = -16'sd53;
gen_input_real[671] = -16'sd57;
gen_input_real[927] = 16'sd51;
gen_input_real[223] = 16'sd59;
gen_input_real[479] = -16'sd43;
gen_input_real[735] = -16'sd46;
gen_input_real[991] = 16'sd33;
gen_input_real[47] = 16'sd27;
gen_input_real[303] = -16'sd17;
gen_input_real[559] = -16'sd15;
gen_input_real[815] = -16'sd3;
gen_input_real[111] = 16'sd10;
gen_input_real[367] = 16'sd15;
gen_input_real[623] = -16'sd17;
gen_input_real[879] = -16'sd8;
gen_input_real[175] = 16'sd32;
gen_input_real[431] = -16'sd5;
gen_input_real[687] = -16'sd37;
gen_input_real[943] = 16'sd11;
gen_input_real[239] = 16'sd26;
gen_input_real[495] = -16'sd4;
gen_input_real[751] = -16'sd20;
gen_input_real[1007] = -16'sd9;
gen_input_real[63] = 16'sd30;
gen_input_real[319] = 16'sd16;
gen_input_real[575] = -16'sd40;
gen_input_real[831] = -16'sd7;
gen_input_real[127] = 16'sd41;
gen_input_real[383] = -16'sd7;
gen_input_real[639] = -16'sd35;
gen_input_real[895] = 16'sd16;
gen_input_real[191] = 16'sd27;
gen_input_real[447] = -16'sd9;
gen_input_real[703] = -16'sd33;
gen_input_real[959] = -16'sd3;
gen_input_real[255] = 16'sd74;
gen_input_real[511] = 16'sd8;
gen_input_real[767] = -16'sd127;
gen_input_real[1023] = 16'sd0;
