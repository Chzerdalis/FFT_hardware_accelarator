0 0
5 -26
34 -83
117 -175
453 -453
-182 122
-170 70
-175 34
-162 0
-175 -34
-170 -70
-182 -122
453 453
117 175
34 83
5 26
