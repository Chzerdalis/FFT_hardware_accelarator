0 0
88 -447
536 -1296
2178 -3260
6904 -6904
-2783 1859
-3060 1267
-2639 525
-2448 0
-2639 -525
-3060 -1267
-2783 -1859
6904 6904
2178 3260
536 1296
88 447
