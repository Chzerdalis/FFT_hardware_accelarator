gen_input_real[0] = 24'sd0;
gen_input_real[16] = 24'sd2047;
gen_input_real[32] = 24'sd123;
gen_input_real[48] = -24'sd1472;
gen_input_real[4] = -24'sd277;
gen_input_real[20] = 24'sd917;
gen_input_real[36] = 24'sd252;
gen_input_real[52] = -24'sd590;
gen_input_real[8] = 24'sd110;
gen_input_real[24] = 24'sd367;
gen_input_real[40] = -24'sd535;
gen_input_real[56] = -24'sd187;
gen_input_real[12] = 24'sd580;
gen_input_real[28] = 24'sd95;
gen_input_real[44] = -24'sd287;
gen_input_real[60] = -24'sd59;
gen_input_real[1] = 24'sd26;
gen_input_real[17] = -24'sd86;
gen_input_real[33] = 24'sd78;
gen_input_real[49] = 24'sd361;
gen_input_real[5] = -24'sd96;
gen_input_real[21] = -24'sd581;
gen_input_real[37] = -24'sd2;
gen_input_real[53] = 24'sd614;
gen_input_real[9] = 24'sd197;
gen_input_real[25] = -24'sd466;
gen_input_real[41] = -24'sd307;
gen_input_real[57] = 24'sd242;
gen_input_real[13] = 24'sd313;
gen_input_real[29] = -24'sd18;
gen_input_real[45] = -24'sd299;
gen_input_real[61] = -24'sd189;
gen_input_real[2] = 24'sd189;
gen_input_real[18] = 24'sd299;
gen_input_real[34] = 24'sd18;
gen_input_real[50] = -24'sd313;
gen_input_real[6] = -24'sd242;
gen_input_real[22] = 24'sd307;
gen_input_real[38] = 24'sd466;
gen_input_real[54] = -24'sd197;
gen_input_real[10] = -24'sd614;
gen_input_real[26] = 24'sd2;
gen_input_real[42] = 24'sd581;
gen_input_real[58] = 24'sd96;
gen_input_real[14] = -24'sd361;
gen_input_real[30] = -24'sd78;
gen_input_real[46] = 24'sd86;
gen_input_real[62] = -24'sd26;
gen_input_real[3] = 24'sd59;
gen_input_real[19] = 24'sd287;
gen_input_real[35] = -24'sd95;
gen_input_real[51] = -24'sd580;
gen_input_real[7] = 24'sd187;
gen_input_real[23] = 24'sd535;
gen_input_real[39] = -24'sd367;
gen_input_real[55] = -24'sd110;
gen_input_real[11] = 24'sd590;
gen_input_real[27] = -24'sd252;
gen_input_real[43] = -24'sd917;
gen_input_real[59] = 24'sd277;
gen_input_real[15] = 24'sd1472;
gen_input_real[31] = -24'sd123;
gen_input_real[47] = -24'sd2047;
gen_input_real[63] = 24'sd0;
