gen_input_real[0] = 32'sd0;
gen_input_real[16] = 32'sd32767;
gen_input_real[32] = 32'sd1981;
gen_input_real[48] = -32'sd23568;
gen_input_real[4] = -32'sd4439;
gen_input_real[20] = 32'sd14684;
gen_input_real[36] = 32'sd4049;
gen_input_real[52] = -32'sd9459;
gen_input_real[8] = 32'sd1765;
gen_input_real[24] = 32'sd5883;
gen_input_real[40] = -32'sd8572;
gen_input_real[56] = -32'sd3008;
gen_input_real[12] = 32'sd9295;
gen_input_real[28] = 32'sd1527;
gen_input_real[44] = -32'sd4595;
gen_input_real[60] = -32'sd960;
gen_input_real[1] = 32'sd423;
gen_input_real[17] = -32'sd1391;
gen_input_real[33] = 32'sd1263;
gen_input_real[49] = 32'sd5791;
gen_input_real[5] = -32'sd1548;
gen_input_real[21] = -32'sd9310;
gen_input_real[37] = -32'sd41;
gen_input_real[53] = 32'sd9838;
gen_input_real[9] = 32'sd3160;
gen_input_real[25] = -32'sd7469;
gen_input_real[41] = -32'sd4922;
gen_input_real[57] = 32'sd3881;
gen_input_real[13] = 32'sd5022;
gen_input_real[29] = -32'sd293;
gen_input_real[45] = -32'sd4797;
gen_input_real[61] = -32'sd3039;
gen_input_real[2] = 32'sd3039;
gen_input_real[18] = 32'sd4797;
gen_input_real[34] = 32'sd293;
gen_input_real[50] = -32'sd5022;
gen_input_real[6] = -32'sd3881;
gen_input_real[22] = 32'sd4922;
gen_input_real[38] = 32'sd7469;
gen_input_real[54] = -32'sd3160;
gen_input_real[10] = -32'sd9838;
gen_input_real[26] = 32'sd41;
gen_input_real[42] = 32'sd9310;
gen_input_real[58] = 32'sd1548;
gen_input_real[14] = -32'sd5791;
gen_input_real[30] = -32'sd1263;
gen_input_real[46] = 32'sd1391;
gen_input_real[62] = -32'sd423;
gen_input_real[3] = 32'sd960;
gen_input_real[19] = 32'sd4595;
gen_input_real[35] = -32'sd1527;
gen_input_real[51] = -32'sd9295;
gen_input_real[7] = 32'sd3008;
gen_input_real[23] = 32'sd8572;
gen_input_real[39] = -32'sd5883;
gen_input_real[55] = -32'sd1765;
gen_input_real[11] = 32'sd9459;
gen_input_real[27] = -32'sd4049;
gen_input_real[43] = -32'sd14684;
gen_input_real[59] = 32'sd4439;
gen_input_real[15] = 32'sd23568;
gen_input_real[31] = -32'sd1981;
gen_input_real[47] = -32'sd32767;
gen_input_real[63] = 32'sd0;
