gen_input_real[0] = 24'sd0;
gen_input_real[256] = 24'sd2047;
gen_input_real[512] = -24'sd130;
gen_input_real[768] = -24'sd1207;
gen_input_real[64] = 24'sd60;
gen_input_real[320] = 24'sd540;
gen_input_real[576] = 24'sd159;
gen_input_real[832] = -24'sd439;
gen_input_real[128] = -24'sd260;
gen_input_real[384] = 24'sd566;
gen_input_real[640] = 24'sd128;
gen_input_real[896] = -24'sd670;
gen_input_real[192] = 24'sd126;
gen_input_real[448] = 24'sd660;
gen_input_real[704] = -24'sd272;
gen_input_real[960] = -24'sd488;
gen_input_real[16] = 24'sd152;
gen_input_real[272] = 24'sd326;
gen_input_real[528] = 24'sd77;
gen_input_real[784] = -24'sd421;
gen_input_real[80] = -24'sd184;
gen_input_real[336] = 24'sd602;
gen_input_real[592] = 24'sd95;
gen_input_real[848] = -24'sd522;
gen_input_real[144] = 24'sd132;
gen_input_real[400] = 24'sd276;
gen_input_real[656] = -24'sd250;
gen_input_real[912] = -24'sd167;
gen_input_real[208] = 24'sd52;
gen_input_real[464] = 24'sd244;
gen_input_real[720] = 24'sd289;
gen_input_real[976] = -24'sd450;
gen_input_real[32] = -24'sd537;
gen_input_real[288] = 24'sd744;
gen_input_real[544] = 24'sd705;
gen_input_real[800] = -24'sd965;
gen_input_real[96] = -24'sd829;
gen_input_real[352] = 24'sd930;
gen_input_real[608] = 24'sd863;
gen_input_real[864] = -24'sd750;
gen_input_real[160] = -24'sd810;
gen_input_real[416] = 24'sd733;
gen_input_real[672] = 24'sd723;
gen_input_real[928] = -24'sd837;
gen_input_real[224] = -24'sd619;
gen_input_real[480] = 24'sd717;
gen_input_real[736] = 24'sd563;
gen_input_real[992] = -24'sd354;
gen_input_real[48] = -24'sd610;
gen_input_real[304] = 24'sd118;
gen_input_real[560] = 24'sd579;
gen_input_real[816] = -24'sd263;
gen_input_real[112] = -24'sd320;
gen_input_real[368] = 24'sd622;
gen_input_real[624] = 24'sd22;
gen_input_real[880] = -24'sd846;
gen_input_real[176] = 24'sd34;
gen_input_real[432] = 24'sd835;
gen_input_real[688] = 24'sd96;
gen_input_real[944] = -24'sd750;
gen_input_real[240] = -24'sd143;
gen_input_real[496] = 24'sd710;
gen_input_real[752] = 24'sd92;
gen_input_real[1008] = -24'sd605;
gen_input_real[4] = -24'sd78;
gen_input_real[260] = 24'sd393;
gen_input_real[516] = 24'sd95;
gen_input_real[772] = -24'sd187;
gen_input_real[68] = -24'sd148;
gen_input_real[324] = 24'sd43;
gen_input_real[580] = 24'sd286;
gen_input_real[836] = -24'sd53;
gen_input_real[132] = -24'sd470;
gen_input_real[388] = 24'sd237;
gen_input_real[644] = 24'sd655;
gen_input_real[900] = -24'sd352;
gen_input_real[196] = -24'sd865;
gen_input_real[452] = 24'sd262;
gen_input_real[708] = 24'sd1028;
gen_input_real[964] = -24'sd77;
gen_input_real[20] = -24'sd938;
gen_input_real[276] = -24'sd142;
gen_input_real[532] = 24'sd654;
gen_input_real[788] = 24'sd391;
gen_input_real[84] = -24'sd445;
gen_input_real[340] = -24'sd522;
gen_input_real[596] = 24'sd309;
gen_input_real[852] = 24'sd338;
gen_input_real[148] = -24'sd258;
gen_input_real[404] = 24'sd86;
gen_input_real[660] = 24'sd486;
gen_input_real[916] = -24'sd447;
gen_input_real[212] = -24'sd788;
gen_input_real[468] = 24'sd611;
gen_input_real[724] = 24'sd778;
gen_input_real[980] = -24'sd643;
gen_input_real[36] = -24'sd546;
gen_input_real[292] = 24'sd598;
gen_input_real[548] = 24'sd400;
gen_input_real[804] = -24'sd515;
gen_input_real[100] = -24'sd422;
gen_input_real[356] = 24'sd429;
gen_input_real[612] = 24'sd483;
gen_input_real[868] = -24'sd430;
gen_input_real[164] = -24'sd430;
gen_input_real[420] = 24'sd473;
gen_input_real[676] = 24'sd225;
gen_input_real[932] = -24'sd325;
gen_input_real[228] = -24'sd53;
gen_input_real[484] = 24'sd34;
gen_input_real[740] = 24'sd232;
gen_input_real[996] = 24'sd142;
gen_input_real[52] = -24'sd634;
gen_input_real[308] = -24'sd164;
gen_input_real[564] = 24'sd700;
gen_input_real[820] = 24'sd111;
gen_input_real[116] = -24'sd296;
gen_input_real[372] = -24'sd69;
gen_input_real[628] = -24'sd143;
gen_input_real[884] = 24'sd153;
gen_input_real[180] = 24'sd273;
gen_input_real[436] = -24'sd379;
gen_input_real[692] = -24'sd175;
gen_input_real[948] = 24'sd563;
gen_input_real[244] = 24'sd53;
gen_input_real[500] = -24'sd540;
gen_input_real[756] = 24'sd64;
gen_input_real[1012] = 24'sd373;
gen_input_real[8] = -24'sd174;
gen_input_real[264] = -24'sd189;
gen_input_real[520] = 24'sd235;
gen_input_real[776] = -24'sd4;
gen_input_real[72] = -24'sd340;
gen_input_real[328] = 24'sd199;
gen_input_real[584] = 24'sd582;
gen_input_real[840] = -24'sd283;
gen_input_real[136] = -24'sd823;
gen_input_real[392] = 24'sd174;
gen_input_real[648] = 24'sd876;
gen_input_real[904] = 24'sd27;
gen_input_real[200] = -24'sd727;
gen_input_real[456] = -24'sd151;
gen_input_real[712] = 24'sd466;
gen_input_real[968] = 24'sd157;
gen_input_real[24] = -24'sd232;
gen_input_real[280] = -24'sd97;
gen_input_real[536] = 24'sd167;
gen_input_real[792] = 24'sd22;
gen_input_real[88] = -24'sd242;
gen_input_real[344] = 24'sd17;
gen_input_real[600] = 24'sd290;
gen_input_real[856] = -24'sd44;
gen_input_real[152] = -24'sd259;
gen_input_real[408] = 24'sd124;
gen_input_real[664] = 24'sd196;
gen_input_real[920] = -24'sd239;
gen_input_real[216] = -24'sd80;
gen_input_real[472] = 24'sd278;
gen_input_real[728] = -24'sd215;
gen_input_real[984] = -24'sd153;
gen_input_real[40] = 24'sd715;
gen_input_real[296] = -24'sd41;
gen_input_real[552] = -24'sd1000;
gen_input_real[808] = 24'sd98;
gen_input_real[104] = 24'sd687;
gen_input_real[360] = 24'sd103;
gen_input_real[616] = -24'sd118;
gen_input_real[872] = -24'sd371;
gen_input_real[168] = -24'sd171;
gen_input_real[424] = 24'sd331;
gen_input_real[680] = 24'sd195;
gen_input_real[936] = -24'sd1;
gen_input_real[232] = -24'sd220;
gen_input_real[488] = -24'sd290;
gen_input_real[744] = 24'sd250;
gen_input_real[1000] = 24'sd441;
gen_input_real[56] = -24'sd193;
gen_input_real[312] = -24'sd418;
gen_input_real[568] = 24'sd125;
gen_input_real[824] = 24'sd229;
gen_input_real[120] = -24'sd31;
gen_input_real[376] = -24'sd134;
gen_input_real[632] = -24'sd122;
gen_input_real[888] = 24'sd277;
gen_input_real[184] = 24'sd117;
gen_input_real[440] = -24'sd423;
gen_input_real[696] = 24'sd88;
gen_input_real[952] = 24'sd335;
gen_input_real[248] = -24'sd240;
gen_input_real[504] = -24'sd64;
gen_input_real[760] = 24'sd265;
gen_input_real[1016] = -24'sd218;
gen_input_real[12] = -24'sd235;
gen_input_real[268] = 24'sd445;
gen_input_real[524] = 24'sd119;
gen_input_real[780] = -24'sd565;
gen_input_real[76] = 24'sd89;
gen_input_real[332] = 24'sd580;
gen_input_real[588] = -24'sd236;
gen_input_real[844] = -24'sd632;
gen_input_real[140] = 24'sd157;
gen_input_real[396] = 24'sd724;
gen_input_real[652] = -24'sd3;
gen_input_real[908] = -24'sd672;
gen_input_real[204] = 24'sd36;
gen_input_real[460] = 24'sd447;
gen_input_real[716] = -24'sd121;
gen_input_real[972] = -24'sd270;
gen_input_real[28] = -24'sd9;
gen_input_real[284] = 24'sd348;
gen_input_real[540] = 24'sd239;
gen_input_real[796] = -24'sd516;
gen_input_real[92] = -24'sd242;
gen_input_real[348] = 24'sd406;
gen_input_real[604] = -24'sd37;
gen_input_real[860] = -24'sd38;
gen_input_real[156] = 24'sd373;
gen_input_real[412] = -24'sd226;
gen_input_real[668] = -24'sd592;
gen_input_real[924] = 24'sd208;
gen_input_real[220] = 24'sd660;
gen_input_real[476] = -24'sd15;
gen_input_real[732] = -24'sd591;
gen_input_real[988] = -24'sd195;
gen_input_real[44] = 24'sd432;
gen_input_real[300] = 24'sd314;
gen_input_real[556] = -24'sd216;
gen_input_real[812] = -24'sd265;
gen_input_real[108] = -24'sd44;
gen_input_real[364] = 24'sd125;
gen_input_real[620] = 24'sd317;
gen_input_real[876] = -24'sd97;
gen_input_real[172] = -24'sd506;
gen_input_real[428] = 24'sd276;
gen_input_real[684] = 24'sd479;
gen_input_real[940] = -24'sd523;
gen_input_real[236] = -24'sd266;
gen_input_real[492] = 24'sd660;
gen_input_real[748] = 24'sd85;
gen_input_real[1004] = -24'sd656;
gen_input_real[60] = -24'sd94;
gen_input_real[316] = 24'sd519;
gen_input_real[572] = 24'sd300;
gen_input_real[828] = -24'sd314;
gen_input_real[124] = -24'sd660;
gen_input_real[380] = 24'sd317;
gen_input_real[636] = 24'sd992;
gen_input_real[892] = -24'sd536;
gen_input_real[188] = -24'sd910;
gen_input_real[444] = 24'sd548;
gen_input_real[700] = 24'sd337;
gen_input_real[956] = -24'sd320;
gen_input_real[252] = 24'sd208;
gen_input_real[508] = 24'sd322;
gen_input_real[764] = -24'sd337;
gen_input_real[1020] = -24'sd646;
gen_input_real[1] = 24'sd206;
gen_input_real[257] = 24'sd907;
gen_input_real[513] = -24'sd102;
gen_input_real[769] = -24'sd948;
gen_input_real[65] = 24'sd149;
gen_input_real[321] = 24'sd896;
gen_input_real[577] = -24'sd260;
gen_input_real[833] = -24'sd711;
gen_input_real[129] = 24'sd236;
gen_input_real[385] = 24'sd425;
gen_input_real[641] = 24'sd1;
gen_input_real[897] = -24'sd315;
gen_input_real[193] = -24'sd378;
gen_input_real[449] = 24'sd399;
gen_input_real[705] = 24'sd648;
gen_input_real[961] = -24'sd486;
gen_input_real[17] = -24'sd568;
gen_input_real[273] = 24'sd543;
gen_input_real[529] = 24'sd284;
gen_input_real[785] = -24'sd471;
gen_input_real[81] = -24'sd165;
gen_input_real[337] = 24'sd163;
gen_input_real[593] = 24'sd310;
gen_input_real[849] = 24'sd148;
gen_input_real[145] = -24'sd521;
gen_input_real[401] = -24'sd165;
gen_input_real[657] = 24'sd654;
gen_input_real[913] = -24'sd33;
gen_input_real[209] = -24'sd718;
gen_input_real[465] = 24'sd128;
gen_input_real[721] = 24'sd687;
gen_input_real[977] = -24'sd81;
gen_input_real[33] = -24'sd622;
gen_input_real[289] = 24'sd152;
gen_input_real[545] = 24'sd695;
gen_input_real[801] = -24'sd378;
gen_input_real[97] = -24'sd760;
gen_input_real[353] = 24'sd573;
gen_input_real[609] = 24'sd568;
gen_input_real[865] = -24'sd706;
gen_input_real[161] = -24'sd299;
gen_input_real[417] = 24'sd851;
gen_input_real[673] = 24'sd271;
gen_input_real[929] = -24'sd989;
gen_input_real[225] = -24'sd494;
gen_input_real[481] = 24'sd1016;
gen_input_real[737] = 24'sd792;
gen_input_real[993] = -24'sd834;
gen_input_real[49] = -24'sd1025;
gen_input_real[305] = 24'sd476;
gen_input_real[561] = 24'sd1073;
gen_input_real[817] = -24'sd189;
gen_input_real[113] = -24'sd882;
gen_input_real[369] = 24'sd189;
gen_input_real[625] = 24'sd586;
gen_input_real[881] = -24'sd343;
gen_input_real[177] = -24'sd392;
gen_input_real[433] = 24'sd381;
gen_input_real[689] = 24'sd307;
gen_input_real[945] = -24'sd301;
gen_input_real[241] = -24'sd211;
gen_input_real[497] = 24'sd215;
gen_input_real[753] = 24'sd155;
gen_input_real[1009] = -24'sd73;
gen_input_real[5] = -24'sd255;
gen_input_real[261] = -24'sd168;
gen_input_real[517] = 24'sd453;
gen_input_real[773] = 24'sd381;
gen_input_real[69] = -24'sd614;
gen_input_real[325] = -24'sd420;
gen_input_real[581] = 24'sd649;
gen_input_real[837] = 24'sd245;
gen_input_real[133] = -24'sd531;
gen_input_real[389] = 24'sd41;
gen_input_real[645] = 24'sd442;
gen_input_real[901] = -24'sd251;
gen_input_real[197] = -24'sd595;
gen_input_real[453] = 24'sd323;
gen_input_real[709] = 24'sd870;
gen_input_real[965] = -24'sd324;
gen_input_real[21] = -24'sd1077;
gen_input_real[277] = 24'sd212;
gen_input_real[533] = 24'sd1242;
gen_input_real[789] = 24'sd25;
gen_input_real[85] = -24'sd1319;
gen_input_real[341] = -24'sd221;
gen_input_real[597] = 24'sd1187;
gen_input_real[853] = 24'sd266;
gen_input_real[149] = -24'sd1011;
gen_input_real[405] = -24'sd197;
gen_input_real[661] = 24'sd1038;
gen_input_real[917] = 24'sd119;
gen_input_real[213] = -24'sd1110;
gen_input_real[469] = -24'sd99;
gen_input_real[725] = 24'sd988;
gen_input_real[981] = 24'sd11;
gen_input_real[37] = -24'sd759;
gen_input_real[293] = 24'sd219;
gen_input_real[549] = 24'sd446;
gen_input_real[805] = -24'sd378;
gen_input_real[101] = -24'sd69;
gen_input_real[357] = 24'sd248;
gen_input_real[613] = 24'sd4;
gen_input_real[869] = 24'sd70;
gen_input_real[165] = -24'sd348;
gen_input_real[421] = -24'sd260;
gen_input_real[677] = 24'sd608;
gen_input_real[933] = 24'sd160;
gen_input_real[229] = -24'sd540;
gen_input_real[485] = 24'sd46;
gen_input_real[741] = 24'sd444;
gen_input_real[997] = -24'sd67;
gen_input_real[53] = -24'sd486;
gen_input_real[309] = -24'sd155;
gen_input_real[565] = 24'sd486;
gen_input_real[821] = 24'sd362;
gen_input_real[117] = -24'sd433;
gen_input_real[373] = -24'sd359;
gen_input_real[629] = 24'sd550;
gen_input_real[885] = 24'sd315;
gen_input_real[181] = -24'sd759;
gen_input_real[437] = -24'sd417;
gen_input_real[693] = 24'sd789;
gen_input_real[949] = 24'sd650;
gen_input_real[245] = -24'sd732;
gen_input_real[501] = -24'sd994;
gen_input_real[757] = 24'sd771;
gen_input_real[1013] = 24'sd1296;
gen_input_real[9] = -24'sd778;
gen_input_real[265] = -24'sd1240;
gen_input_real[521] = 24'sd643;
gen_input_real[777] = 24'sd800;
gen_input_real[73] = -24'sd504;
gen_input_real[329] = -24'sd286;
gen_input_real[585] = 24'sd460;
gen_input_real[841] = -24'sd48;
gen_input_real[137] = -24'sd465;
gen_input_real[393] = 24'sd143;
gen_input_real[649] = 24'sd540;
gen_input_real[905] = -24'sd21;
gen_input_real[201] = -24'sd672;
gen_input_real[457] = -24'sd207;
gen_input_real[713] = 24'sd666;
gen_input_real[969] = 24'sd342;
gen_input_real[25] = -24'sd518;
gen_input_real[281] = -24'sd317;
gen_input_real[537] = 24'sd505;
gen_input_real[793] = 24'sd262;
gen_input_real[89] = -24'sd656;
gen_input_real[345] = -24'sd194;
gen_input_real[601] = 24'sd644;
gen_input_real[857] = 24'sd9;
gen_input_real[153] = -24'sd368;
gen_input_real[409] = 24'sd110;
gen_input_real[665] = 24'sd157;
gen_input_real[921] = 24'sd128;
gen_input_real[217] = -24'sd258;
gen_input_real[473] = -24'sd527;
gen_input_real[729] = 24'sd429;
gen_input_real[985] = 24'sd719;
gen_input_real[41] = -24'sd250;
gen_input_real[297] = -24'sd770;
gen_input_real[553] = -24'sd215;
gen_input_real[809] = 24'sd854;
gen_input_real[105] = 24'sd501;
gen_input_real[361] = -24'sd899;
gen_input_real[617] = -24'sd427;
gen_input_real[873] = 24'sd864;
gen_input_real[169] = 24'sd137;
gen_input_real[425] = -24'sd805;
gen_input_real[681] = 24'sd195;
gen_input_real[937] = 24'sd602;
gen_input_real[233] = -24'sd331;
gen_input_real[489] = -24'sd253;
gen_input_real[745] = 24'sd162;
gen_input_real[1001] = 24'sd116;
gen_input_real[57] = 24'sd26;
gen_input_real[313] = -24'sd325;
gen_input_real[569] = 24'sd70;
gen_input_real[825] = 24'sd562;
gen_input_real[121] = -24'sd388;
gen_input_real[377] = -24'sd642;
gen_input_real[633] = 24'sd677;
gen_input_real[889] = 24'sd651;
gen_input_real[185] = -24'sd762;
gen_input_real[441] = -24'sd603;
gen_input_real[697] = 24'sd620;
gen_input_real[953] = 24'sd550;
gen_input_real[249] = -24'sd377;
gen_input_real[505] = -24'sd544;
gen_input_real[761] = 24'sd269;
gen_input_real[1017] = 24'sd448;
gen_input_real[13] = -24'sd372;
gen_input_real[269] = -24'sd203;
gen_input_real[525] = 24'sd397;
gen_input_real[781] = -24'sd16;
gen_input_real[77] = -24'sd88;
gen_input_real[333] = 24'sd14;
gen_input_real[589] = -24'sd334;
gen_input_real[845] = 24'sd198;
gen_input_real[141] = 24'sd432;
gen_input_real[397] = -24'sd398;
gen_input_real[653] = -24'sd206;
gen_input_real[909] = 24'sd412;
gen_input_real[205] = 24'sd161;
gen_input_real[461] = -24'sd254;
gen_input_real[717] = -24'sd474;
gen_input_real[973] = 24'sd41;
gen_input_real[29] = 24'sd679;
gen_input_real[285] = 24'sd112;
gen_input_real[541] = -24'sd451;
gen_input_real[797] = -24'sd175;
gen_input_real[93] = 24'sd15;
gen_input_real[349] = 24'sd161;
gen_input_real[605] = 24'sd277;
gen_input_real[861] = -24'sd18;
gen_input_real[157] = -24'sd240;
gen_input_real[413] = -24'sd295;
gen_input_real[669] = -24'sd79;
gen_input_real[925] = 24'sd678;
gen_input_real[221] = 24'sd361;
gen_input_real[477] = -24'sd968;
gen_input_real[733] = -24'sd317;
gen_input_real[989] = 24'sd1043;
gen_input_real[45] = 24'sd26;
gen_input_real[301] = -24'sd849;
gen_input_real[557] = 24'sd193;
gen_input_real[813] = 24'sd469;
gen_input_real[109] = -24'sd187;
gen_input_real[365] = -24'sd157;
gen_input_real[621] = 24'sd99;
gen_input_real[877] = 24'sd142;
gen_input_real[173] = -24'sd44;
gen_input_real[429] = -24'sd304;
gen_input_real[685] = 24'sd9;
gen_input_real[941] = 24'sd339;
gen_input_real[237] = -24'sd42;
gen_input_real[493] = -24'sd167;
gen_input_real[749] = 24'sd108;
gen_input_real[1005] = -24'sd87;
gen_input_real[61] = 24'sd4;
gen_input_real[317] = 24'sd267;
gen_input_real[573] = -24'sd231;
gen_input_real[829] = -24'sd297;
gen_input_real[125] = 24'sd163;
gen_input_real[381] = 24'sd281;
gen_input_real[637] = 24'sd263;
gen_input_real[893] = -24'sd326;
gen_input_real[189] = -24'sd596;
gen_input_real[445] = 24'sd351;
gen_input_real[701] = 24'sd539;
gen_input_real[957] = -24'sd325;
gen_input_real[253] = -24'sd241;
gen_input_real[509] = 24'sd320;
gen_input_real[765] = -24'sd61;
gen_input_real[1021] = -24'sd261;
gen_input_real[2] = 24'sd261;
gen_input_real[258] = 24'sd61;
gen_input_real[514] = -24'sd320;
gen_input_real[770] = 24'sd241;
gen_input_real[66] = 24'sd325;
gen_input_real[322] = -24'sd539;
gen_input_real[578] = -24'sd351;
gen_input_real[834] = 24'sd596;
gen_input_real[130] = 24'sd326;
gen_input_real[386] = -24'sd263;
gen_input_real[642] = -24'sd281;
gen_input_real[898] = -24'sd163;
gen_input_real[194] = 24'sd297;
gen_input_real[450] = 24'sd231;
gen_input_real[706] = -24'sd267;
gen_input_real[962] = -24'sd4;
gen_input_real[18] = 24'sd87;
gen_input_real[274] = -24'sd108;
gen_input_real[530] = 24'sd167;
gen_input_real[786] = 24'sd42;
gen_input_real[82] = -24'sd339;
gen_input_real[338] = -24'sd9;
gen_input_real[594] = 24'sd304;
gen_input_real[850] = 24'sd44;
gen_input_real[146] = -24'sd142;
gen_input_real[402] = -24'sd99;
gen_input_real[658] = 24'sd157;
gen_input_real[914] = 24'sd187;
gen_input_real[210] = -24'sd469;
gen_input_real[466] = -24'sd193;
gen_input_real[722] = 24'sd849;
gen_input_real[978] = -24'sd26;
gen_input_real[34] = -24'sd1043;
gen_input_real[290] = 24'sd317;
gen_input_real[546] = 24'sd968;
gen_input_real[802] = -24'sd361;
gen_input_real[98] = -24'sd678;
gen_input_real[354] = 24'sd79;
gen_input_real[610] = 24'sd295;
gen_input_real[866] = 24'sd240;
gen_input_real[162] = 24'sd18;
gen_input_real[418] = -24'sd277;
gen_input_real[674] = -24'sd161;
gen_input_real[930] = -24'sd15;
gen_input_real[226] = 24'sd175;
gen_input_real[482] = 24'sd451;
gen_input_real[738] = -24'sd112;
gen_input_real[994] = -24'sd679;
gen_input_real[50] = -24'sd41;
gen_input_real[306] = 24'sd474;
gen_input_real[562] = 24'sd254;
gen_input_real[818] = -24'sd161;
gen_input_real[114] = -24'sd412;
gen_input_real[370] = 24'sd206;
gen_input_real[626] = 24'sd398;
gen_input_real[882] = -24'sd432;
gen_input_real[178] = -24'sd198;
gen_input_real[434] = 24'sd334;
gen_input_real[690] = -24'sd14;
gen_input_real[946] = 24'sd88;
gen_input_real[242] = 24'sd16;
gen_input_real[498] = -24'sd397;
gen_input_real[754] = 24'sd203;
gen_input_real[1010] = 24'sd372;
gen_input_real[6] = -24'sd448;
gen_input_real[262] = -24'sd269;
gen_input_real[518] = 24'sd544;
gen_input_real[774] = 24'sd377;
gen_input_real[70] = -24'sd550;
gen_input_real[326] = -24'sd620;
gen_input_real[582] = 24'sd603;
gen_input_real[838] = 24'sd762;
gen_input_real[134] = -24'sd651;
gen_input_real[390] = -24'sd677;
gen_input_real[646] = 24'sd642;
gen_input_real[902] = 24'sd388;
gen_input_real[198] = -24'sd562;
gen_input_real[454] = -24'sd70;
gen_input_real[710] = 24'sd325;
gen_input_real[966] = -24'sd26;
gen_input_real[22] = -24'sd116;
gen_input_real[278] = -24'sd162;
gen_input_real[534] = 24'sd253;
gen_input_real[790] = 24'sd331;
gen_input_real[86] = -24'sd602;
gen_input_real[342] = -24'sd195;
gen_input_real[598] = 24'sd805;
gen_input_real[854] = -24'sd137;
gen_input_real[150] = -24'sd864;
gen_input_real[406] = 24'sd427;
gen_input_real[662] = 24'sd899;
gen_input_real[918] = -24'sd501;
gen_input_real[214] = -24'sd854;
gen_input_real[470] = 24'sd215;
gen_input_real[726] = 24'sd770;
gen_input_real[982] = 24'sd250;
gen_input_real[38] = -24'sd719;
gen_input_real[294] = -24'sd429;
gen_input_real[550] = 24'sd527;
gen_input_real[806] = 24'sd258;
gen_input_real[102] = -24'sd128;
gen_input_real[358] = -24'sd157;
gen_input_real[614] = -24'sd110;
gen_input_real[870] = 24'sd368;
gen_input_real[166] = -24'sd9;
gen_input_real[422] = -24'sd644;
gen_input_real[678] = 24'sd194;
gen_input_real[934] = 24'sd656;
gen_input_real[230] = -24'sd262;
gen_input_real[486] = -24'sd505;
gen_input_real[742] = 24'sd317;
gen_input_real[998] = 24'sd518;
gen_input_real[54] = -24'sd342;
gen_input_real[310] = -24'sd666;
gen_input_real[566] = 24'sd207;
gen_input_real[822] = 24'sd672;
gen_input_real[118] = 24'sd21;
gen_input_real[374] = -24'sd540;
gen_input_real[630] = -24'sd143;
gen_input_real[886] = 24'sd465;
gen_input_real[182] = 24'sd48;
gen_input_real[438] = -24'sd460;
gen_input_real[694] = 24'sd286;
gen_input_real[950] = 24'sd504;
gen_input_real[246] = -24'sd800;
gen_input_real[502] = -24'sd643;
gen_input_real[758] = 24'sd1240;
gen_input_real[1014] = 24'sd778;
gen_input_real[10] = -24'sd1296;
gen_input_real[266] = -24'sd771;
gen_input_real[522] = 24'sd994;
gen_input_real[778] = 24'sd732;
gen_input_real[74] = -24'sd650;
gen_input_real[330] = -24'sd789;
gen_input_real[586] = 24'sd417;
gen_input_real[842] = 24'sd759;
gen_input_real[138] = -24'sd315;
gen_input_real[394] = -24'sd550;
gen_input_real[650] = 24'sd359;
gen_input_real[906] = 24'sd433;
gen_input_real[202] = -24'sd362;
gen_input_real[458] = -24'sd486;
gen_input_real[714] = 24'sd155;
gen_input_real[970] = 24'sd486;
gen_input_real[26] = 24'sd67;
gen_input_real[282] = -24'sd444;
gen_input_real[538] = -24'sd46;
gen_input_real[794] = 24'sd540;
gen_input_real[90] = -24'sd160;
gen_input_real[346] = -24'sd608;
gen_input_real[602] = 24'sd260;
gen_input_real[858] = 24'sd348;
gen_input_real[154] = -24'sd70;
gen_input_real[410] = -24'sd4;
gen_input_real[666] = -24'sd248;
gen_input_real[922] = 24'sd69;
gen_input_real[218] = 24'sd378;
gen_input_real[474] = -24'sd446;
gen_input_real[730] = -24'sd219;
gen_input_real[986] = 24'sd759;
gen_input_real[42] = -24'sd11;
gen_input_real[298] = -24'sd988;
gen_input_real[554] = 24'sd99;
gen_input_real[810] = 24'sd1110;
gen_input_real[106] = -24'sd119;
gen_input_real[362] = -24'sd1038;
gen_input_real[618] = 24'sd197;
gen_input_real[874] = 24'sd1011;
gen_input_real[170] = -24'sd266;
gen_input_real[426] = -24'sd1187;
gen_input_real[682] = 24'sd221;
gen_input_real[938] = 24'sd1319;
gen_input_real[234] = -24'sd25;
gen_input_real[490] = -24'sd1242;
gen_input_real[746] = -24'sd212;
gen_input_real[1002] = 24'sd1077;
gen_input_real[58] = 24'sd324;
gen_input_real[314] = -24'sd870;
gen_input_real[570] = -24'sd323;
gen_input_real[826] = 24'sd595;
gen_input_real[122] = 24'sd251;
gen_input_real[378] = -24'sd442;
gen_input_real[634] = -24'sd41;
gen_input_real[890] = 24'sd531;
gen_input_real[186] = -24'sd245;
gen_input_real[442] = -24'sd649;
gen_input_real[698] = 24'sd420;
gen_input_real[954] = 24'sd614;
gen_input_real[250] = -24'sd381;
gen_input_real[506] = -24'sd453;
gen_input_real[762] = 24'sd168;
gen_input_real[1018] = 24'sd255;
gen_input_real[14] = 24'sd73;
gen_input_real[270] = -24'sd155;
gen_input_real[526] = -24'sd215;
gen_input_real[782] = 24'sd211;
gen_input_real[78] = 24'sd301;
gen_input_real[334] = -24'sd307;
gen_input_real[590] = -24'sd381;
gen_input_real[846] = 24'sd392;
gen_input_real[142] = 24'sd343;
gen_input_real[398] = -24'sd586;
gen_input_real[654] = -24'sd189;
gen_input_real[910] = 24'sd882;
gen_input_real[206] = 24'sd189;
gen_input_real[462] = -24'sd1073;
gen_input_real[718] = -24'sd476;
gen_input_real[974] = 24'sd1025;
gen_input_real[30] = 24'sd834;
gen_input_real[286] = -24'sd792;
gen_input_real[542] = -24'sd1016;
gen_input_real[798] = 24'sd494;
gen_input_real[94] = 24'sd989;
gen_input_real[350] = -24'sd271;
gen_input_real[606] = -24'sd851;
gen_input_real[862] = 24'sd299;
gen_input_real[158] = 24'sd706;
gen_input_real[414] = -24'sd568;
gen_input_real[670] = -24'sd573;
gen_input_real[926] = 24'sd760;
gen_input_real[222] = 24'sd378;
gen_input_real[478] = -24'sd695;
gen_input_real[734] = -24'sd152;
gen_input_real[990] = 24'sd622;
gen_input_real[46] = 24'sd81;
gen_input_real[302] = -24'sd687;
gen_input_real[558] = -24'sd128;
gen_input_real[814] = 24'sd718;
gen_input_real[110] = 24'sd33;
gen_input_real[366] = -24'sd654;
gen_input_real[622] = 24'sd165;
gen_input_real[878] = 24'sd521;
gen_input_real[174] = -24'sd148;
gen_input_real[430] = -24'sd310;
gen_input_real[686] = -24'sd163;
gen_input_real[942] = 24'sd165;
gen_input_real[238] = 24'sd471;
gen_input_real[494] = -24'sd284;
gen_input_real[750] = -24'sd543;
gen_input_real[1006] = 24'sd568;
gen_input_real[62] = 24'sd486;
gen_input_real[318] = -24'sd648;
gen_input_real[574] = -24'sd399;
gen_input_real[830] = 24'sd378;
gen_input_real[126] = 24'sd315;
gen_input_real[382] = -24'sd1;
gen_input_real[638] = -24'sd425;
gen_input_real[894] = -24'sd236;
gen_input_real[190] = 24'sd711;
gen_input_real[446] = 24'sd260;
gen_input_real[702] = -24'sd896;
gen_input_real[958] = -24'sd149;
gen_input_real[254] = 24'sd948;
gen_input_real[510] = 24'sd102;
gen_input_real[766] = -24'sd907;
gen_input_real[1022] = -24'sd206;
gen_input_real[3] = 24'sd646;
gen_input_real[259] = 24'sd337;
gen_input_real[515] = -24'sd322;
gen_input_real[771] = -24'sd208;
gen_input_real[67] = 24'sd320;
gen_input_real[323] = -24'sd337;
gen_input_real[579] = -24'sd548;
gen_input_real[835] = 24'sd910;
gen_input_real[131] = 24'sd536;
gen_input_real[387] = -24'sd992;
gen_input_real[643] = -24'sd317;
gen_input_real[899] = 24'sd660;
gen_input_real[195] = 24'sd314;
gen_input_real[451] = -24'sd300;
gen_input_real[707] = -24'sd519;
gen_input_real[963] = 24'sd94;
gen_input_real[19] = 24'sd656;
gen_input_real[275] = -24'sd85;
gen_input_real[531] = -24'sd660;
gen_input_real[787] = 24'sd266;
gen_input_real[83] = 24'sd523;
gen_input_real[339] = -24'sd479;
gen_input_real[595] = -24'sd276;
gen_input_real[851] = 24'sd506;
gen_input_real[147] = 24'sd97;
gen_input_real[403] = -24'sd317;
gen_input_real[659] = -24'sd125;
gen_input_real[915] = 24'sd44;
gen_input_real[211] = 24'sd265;
gen_input_real[467] = 24'sd216;
gen_input_real[723] = -24'sd314;
gen_input_real[979] = -24'sd432;
gen_input_real[35] = 24'sd195;
gen_input_real[291] = 24'sd591;
gen_input_real[547] = 24'sd15;
gen_input_real[803] = -24'sd660;
gen_input_real[99] = -24'sd208;
gen_input_real[355] = 24'sd592;
gen_input_real[611] = 24'sd226;
gen_input_real[867] = -24'sd373;
gen_input_real[163] = 24'sd38;
gen_input_real[419] = 24'sd37;
gen_input_real[675] = -24'sd406;
gen_input_real[931] = 24'sd242;
gen_input_real[227] = 24'sd516;
gen_input_real[483] = -24'sd239;
gen_input_real[739] = -24'sd348;
gen_input_real[995] = 24'sd9;
gen_input_real[51] = 24'sd270;
gen_input_real[307] = 24'sd121;
gen_input_real[563] = -24'sd447;
gen_input_real[819] = -24'sd36;
gen_input_real[115] = 24'sd672;
gen_input_real[371] = 24'sd3;
gen_input_real[627] = -24'sd724;
gen_input_real[883] = -24'sd157;
gen_input_real[179] = 24'sd632;
gen_input_real[435] = 24'sd236;
gen_input_real[691] = -24'sd580;
gen_input_real[947] = -24'sd89;
gen_input_real[243] = 24'sd565;
gen_input_real[499] = -24'sd119;
gen_input_real[755] = -24'sd445;
gen_input_real[1011] = 24'sd235;
gen_input_real[7] = 24'sd218;
gen_input_real[263] = -24'sd265;
gen_input_real[519] = 24'sd64;
gen_input_real[775] = 24'sd240;
gen_input_real[71] = -24'sd335;
gen_input_real[327] = -24'sd88;
gen_input_real[583] = 24'sd423;
gen_input_real[839] = -24'sd117;
gen_input_real[135] = -24'sd277;
gen_input_real[391] = 24'sd122;
gen_input_real[647] = 24'sd134;
gen_input_real[903] = 24'sd31;
gen_input_real[199] = -24'sd229;
gen_input_real[455] = -24'sd125;
gen_input_real[711] = 24'sd418;
gen_input_real[967] = 24'sd193;
gen_input_real[23] = -24'sd441;
gen_input_real[279] = -24'sd250;
gen_input_real[535] = 24'sd290;
gen_input_real[791] = 24'sd220;
gen_input_real[87] = 24'sd1;
gen_input_real[343] = -24'sd195;
gen_input_real[599] = -24'sd331;
gen_input_real[855] = 24'sd171;
gen_input_real[151] = 24'sd371;
gen_input_real[407] = 24'sd118;
gen_input_real[663] = -24'sd103;
gen_input_real[919] = -24'sd687;
gen_input_real[215] = -24'sd98;
gen_input_real[471] = 24'sd1000;
gen_input_real[727] = 24'sd41;
gen_input_real[983] = -24'sd715;
gen_input_real[39] = 24'sd153;
gen_input_real[295] = 24'sd215;
gen_input_real[551] = -24'sd278;
gen_input_real[807] = 24'sd80;
gen_input_real[103] = 24'sd239;
gen_input_real[359] = -24'sd196;
gen_input_real[615] = -24'sd124;
gen_input_real[871] = 24'sd259;
gen_input_real[167] = 24'sd44;
gen_input_real[423] = -24'sd290;
gen_input_real[679] = -24'sd17;
gen_input_real[935] = 24'sd242;
gen_input_real[231] = -24'sd22;
gen_input_real[487] = -24'sd167;
gen_input_real[743] = 24'sd97;
gen_input_real[999] = 24'sd232;
gen_input_real[55] = -24'sd157;
gen_input_real[311] = -24'sd466;
gen_input_real[567] = 24'sd151;
gen_input_real[823] = 24'sd727;
gen_input_real[119] = -24'sd27;
gen_input_real[375] = -24'sd876;
gen_input_real[631] = -24'sd174;
gen_input_real[887] = 24'sd823;
gen_input_real[183] = 24'sd283;
gen_input_real[439] = -24'sd582;
gen_input_real[695] = -24'sd199;
gen_input_real[951] = 24'sd340;
gen_input_real[247] = 24'sd4;
gen_input_real[503] = -24'sd235;
gen_input_real[759] = 24'sd189;
gen_input_real[1015] = 24'sd174;
gen_input_real[11] = -24'sd373;
gen_input_real[267] = -24'sd64;
gen_input_real[523] = 24'sd540;
gen_input_real[779] = -24'sd53;
gen_input_real[75] = -24'sd563;
gen_input_real[331] = 24'sd175;
gen_input_real[587] = 24'sd379;
gen_input_real[843] = -24'sd273;
gen_input_real[139] = -24'sd153;
gen_input_real[395] = 24'sd143;
gen_input_real[651] = 24'sd69;
gen_input_real[907] = 24'sd296;
gen_input_real[203] = -24'sd111;
gen_input_real[459] = -24'sd700;
gen_input_real[715] = 24'sd164;
gen_input_real[971] = 24'sd634;
gen_input_real[27] = -24'sd142;
gen_input_real[283] = -24'sd232;
gen_input_real[539] = -24'sd34;
gen_input_real[795] = 24'sd53;
gen_input_real[91] = 24'sd325;
gen_input_real[347] = -24'sd225;
gen_input_real[603] = -24'sd473;
gen_input_real[859] = 24'sd430;
gen_input_real[155] = 24'sd430;
gen_input_real[411] = -24'sd483;
gen_input_real[667] = -24'sd429;
gen_input_real[923] = 24'sd422;
gen_input_real[219] = 24'sd515;
gen_input_real[475] = -24'sd400;
gen_input_real[731] = -24'sd598;
gen_input_real[987] = 24'sd546;
gen_input_real[43] = 24'sd643;
gen_input_real[299] = -24'sd778;
gen_input_real[555] = -24'sd611;
gen_input_real[811] = 24'sd788;
gen_input_real[107] = 24'sd447;
gen_input_real[363] = -24'sd486;
gen_input_real[619] = -24'sd86;
gen_input_real[875] = 24'sd258;
gen_input_real[171] = -24'sd338;
gen_input_real[427] = -24'sd309;
gen_input_real[683] = 24'sd522;
gen_input_real[939] = 24'sd445;
gen_input_real[235] = -24'sd391;
gen_input_real[491] = -24'sd654;
gen_input_real[747] = 24'sd142;
gen_input_real[1003] = 24'sd938;
gen_input_real[59] = 24'sd77;
gen_input_real[315] = -24'sd1028;
gen_input_real[571] = -24'sd262;
gen_input_real[827] = 24'sd865;
gen_input_real[123] = 24'sd352;
gen_input_real[379] = -24'sd655;
gen_input_real[635] = -24'sd237;
gen_input_real[891] = 24'sd470;
gen_input_real[187] = 24'sd53;
gen_input_real[443] = -24'sd286;
gen_input_real[699] = -24'sd43;
gen_input_real[955] = 24'sd148;
gen_input_real[251] = 24'sd187;
gen_input_real[507] = -24'sd95;
gen_input_real[763] = -24'sd393;
gen_input_real[1019] = 24'sd78;
gen_input_real[15] = 24'sd605;
gen_input_real[271] = -24'sd92;
gen_input_real[527] = -24'sd710;
gen_input_real[783] = 24'sd143;
gen_input_real[79] = 24'sd750;
gen_input_real[335] = -24'sd96;
gen_input_real[591] = -24'sd835;
gen_input_real[847] = -24'sd34;
gen_input_real[143] = 24'sd846;
gen_input_real[399] = -24'sd22;
gen_input_real[655] = -24'sd622;
gen_input_real[911] = 24'sd320;
gen_input_real[207] = 24'sd263;
gen_input_real[463] = -24'sd579;
gen_input_real[719] = -24'sd118;
gen_input_real[975] = 24'sd610;
gen_input_real[31] = 24'sd354;
gen_input_real[287] = -24'sd563;
gen_input_real[543] = -24'sd717;
gen_input_real[799] = 24'sd619;
gen_input_real[95] = 24'sd837;
gen_input_real[351] = -24'sd723;
gen_input_real[607] = -24'sd733;
gen_input_real[863] = 24'sd810;
gen_input_real[159] = 24'sd750;
gen_input_real[415] = -24'sd863;
gen_input_real[671] = -24'sd930;
gen_input_real[927] = 24'sd829;
gen_input_real[223] = 24'sd965;
gen_input_real[479] = -24'sd705;
gen_input_real[735] = -24'sd744;
gen_input_real[991] = 24'sd537;
gen_input_real[47] = 24'sd450;
gen_input_real[303] = -24'sd289;
gen_input_real[559] = -24'sd244;
gen_input_real[815] = -24'sd52;
gen_input_real[111] = 24'sd167;
gen_input_real[367] = 24'sd250;
gen_input_real[623] = -24'sd276;
gen_input_real[879] = -24'sd132;
gen_input_real[175] = 24'sd522;
gen_input_real[431] = -24'sd95;
gen_input_real[687] = -24'sd602;
gen_input_real[943] = 24'sd184;
gen_input_real[239] = 24'sd421;
gen_input_real[495] = -24'sd77;
gen_input_real[751] = -24'sd326;
gen_input_real[1007] = -24'sd152;
gen_input_real[63] = 24'sd488;
gen_input_real[319] = 24'sd272;
gen_input_real[575] = -24'sd660;
gen_input_real[831] = -24'sd126;
gen_input_real[127] = 24'sd670;
gen_input_real[383] = -24'sd128;
gen_input_real[639] = -24'sd566;
gen_input_real[895] = 24'sd260;
gen_input_real[191] = 24'sd439;
gen_input_real[447] = -24'sd159;
gen_input_real[703] = -24'sd540;
gen_input_real[959] = -24'sd60;
gen_input_real[255] = 24'sd1207;
gen_input_real[511] = 24'sd130;
gen_input_real[767] = -24'sd2047;
gen_input_real[1023] = 24'sd0;
