w_real[0] = 12'h7FF; w_imag[0] = 12'h000;
w_real[1] = 12'h7FF; w_imag[1] = 12'hFCE;
w_real[2] = 12'h7FD; w_imag[2] = 12'hF9C;
w_real[3] = 12'h7FA; w_imag[3] = 12'hF6A;
w_real[4] = 12'h7F6; w_imag[4] = 12'hF38;
w_real[5] = 12'h7F0; w_imag[5] = 12'hF06;
w_real[6] = 12'h7E9; w_imag[6] = 12'hED4;
w_real[7] = 12'h7E1; w_imag[7] = 12'hEA2;
w_real[8] = 12'h7D8; w_imag[8] = 12'hE71;
w_real[9] = 12'h7CE; w_imag[9] = 12'hE40;
w_real[10] = 12'h7C2; w_imag[10] = 12'hE0F;
w_real[11] = 12'h7B5; w_imag[11] = 12'hDDE;
w_real[12] = 12'h7A7; w_imag[12] = 12'hDAE;
w_real[13] = 12'h798; w_imag[13] = 12'hD7E;
w_real[14] = 12'h788; w_imag[14] = 12'hD4F;
w_real[15] = 12'h776; w_imag[15] = 12'hD1F;
w_real[16] = 12'h764; w_imag[16] = 12'hCF1;
w_real[17] = 12'h750; w_imag[17] = 12'hCC3;
w_real[18] = 12'h73B; w_imag[18] = 12'hC95;
w_real[19] = 12'h725; w_imag[19] = 12'hC68;
w_real[20] = 12'h70E; w_imag[20] = 12'hC3B;
w_real[21] = 12'h6F5; w_imag[21] = 12'hC0F;
w_real[22] = 12'h6DC; w_imag[22] = 12'hBE4;
w_real[23] = 12'h6C2; w_imag[23] = 12'hBB9;
w_real[24] = 12'h6A6; w_imag[24] = 12'hB8F;
w_real[25] = 12'h68A; w_imag[25] = 12'hB65;
w_real[26] = 12'h66C; w_imag[26] = 12'hB3D;
w_real[27] = 12'h64E; w_imag[27] = 12'hB15;
w_real[28] = 12'h62F; w_imag[28] = 12'hAED;
w_real[29] = 12'h60E; w_imag[29] = 12'hAC7;
w_real[30] = 12'h5ED; w_imag[30] = 12'hAA1;
w_real[31] = 12'h5CB; w_imag[31] = 12'hA7C;
w_real[32] = 12'h5A8; w_imag[32] = 12'hA58;
w_real[33] = 12'h584; w_imag[33] = 12'hA35;
w_real[34] = 12'h55F; w_imag[34] = 12'hA13;
w_real[35] = 12'h539; w_imag[35] = 12'h9F2;
w_real[36] = 12'h513; w_imag[36] = 12'h9D1;
w_real[37] = 12'h4EB; w_imag[37] = 12'h9B2;
w_real[38] = 12'h4C3; w_imag[38] = 12'h994;
w_real[39] = 12'h49B; w_imag[39] = 12'h976;
w_real[40] = 12'h471; w_imag[40] = 12'h95A;
w_real[41] = 12'h447; w_imag[41] = 12'h93E;
w_real[42] = 12'h41C; w_imag[42] = 12'h924;
w_real[43] = 12'h3F1; w_imag[43] = 12'h90B;
w_real[44] = 12'h3C5; w_imag[44] = 12'h8F2;
w_real[45] = 12'h398; w_imag[45] = 12'h8DB;
w_real[46] = 12'h36B; w_imag[46] = 12'h8C5;
w_real[47] = 12'h33D; w_imag[47] = 12'h8B0;
w_real[48] = 12'h30F; w_imag[48] = 12'h89C;
w_real[49] = 12'h2E1; w_imag[49] = 12'h88A;
w_real[50] = 12'h2B1; w_imag[50] = 12'h878;
w_real[51] = 12'h282; w_imag[51] = 12'h868;
w_real[52] = 12'h252; w_imag[52] = 12'h859;
w_real[53] = 12'h222; w_imag[53] = 12'h84B;
w_real[54] = 12'h1F1; w_imag[54] = 12'h83E;
w_real[55] = 12'h1C0; w_imag[55] = 12'h832;
w_real[56] = 12'h18F; w_imag[56] = 12'h828;
w_real[57] = 12'h15E; w_imag[57] = 12'h81F;
w_real[58] = 12'h12C; w_imag[58] = 12'h817;
w_real[59] = 12'h0FA; w_imag[59] = 12'h810;
w_real[60] = 12'h0C8; w_imag[60] = 12'h80A;
w_real[61] = 12'h096; w_imag[61] = 12'h806;
w_real[62] = 12'h064; w_imag[62] = 12'h803;
w_real[63] = 12'h032; w_imag[63] = 12'h801;
w_real[64] = 12'h000; w_imag[64] = 12'h800;
w_real[65] = 12'hFCE; w_imag[65] = 12'h801;
w_real[66] = 12'hF9C; w_imag[66] = 12'h803;
w_real[67] = 12'hF6A; w_imag[67] = 12'h806;
w_real[68] = 12'hF38; w_imag[68] = 12'h80A;
w_real[69] = 12'hF06; w_imag[69] = 12'h810;
w_real[70] = 12'hED4; w_imag[70] = 12'h817;
w_real[71] = 12'hEA2; w_imag[71] = 12'h81F;
w_real[72] = 12'hE71; w_imag[72] = 12'h828;
w_real[73] = 12'hE40; w_imag[73] = 12'h832;
w_real[74] = 12'hE0F; w_imag[74] = 12'h83E;
w_real[75] = 12'hDDE; w_imag[75] = 12'h84B;
w_real[76] = 12'hDAE; w_imag[76] = 12'h859;
w_real[77] = 12'hD7E; w_imag[77] = 12'h868;
w_real[78] = 12'hD4F; w_imag[78] = 12'h878;
w_real[79] = 12'hD1F; w_imag[79] = 12'h88A;
w_real[80] = 12'hCF1; w_imag[80] = 12'h89C;
w_real[81] = 12'hCC3; w_imag[81] = 12'h8B0;
w_real[82] = 12'hC95; w_imag[82] = 12'h8C5;
w_real[83] = 12'hC68; w_imag[83] = 12'h8DB;
w_real[84] = 12'hC3B; w_imag[84] = 12'h8F2;
w_real[85] = 12'hC0F; w_imag[85] = 12'h90B;
w_real[86] = 12'hBE4; w_imag[86] = 12'h924;
w_real[87] = 12'hBB9; w_imag[87] = 12'h93E;
w_real[88] = 12'hB8F; w_imag[88] = 12'h95A;
w_real[89] = 12'hB65; w_imag[89] = 12'h976;
w_real[90] = 12'hB3D; w_imag[90] = 12'h994;
w_real[91] = 12'hB15; w_imag[91] = 12'h9B2;
w_real[92] = 12'hAED; w_imag[92] = 12'h9D1;
w_real[93] = 12'hAC7; w_imag[93] = 12'h9F2;
w_real[94] = 12'hAA1; w_imag[94] = 12'hA13;
w_real[95] = 12'hA7C; w_imag[95] = 12'hA35;
w_real[96] = 12'hA58; w_imag[96] = 12'hA58;
w_real[97] = 12'hA35; w_imag[97] = 12'hA7C;
w_real[98] = 12'hA13; w_imag[98] = 12'hAA1;
w_real[99] = 12'h9F2; w_imag[99] = 12'hAC7;
w_real[100] = 12'h9D1; w_imag[100] = 12'hAED;
w_real[101] = 12'h9B2; w_imag[101] = 12'hB15;
w_real[102] = 12'h994; w_imag[102] = 12'hB3D;
w_real[103] = 12'h976; w_imag[103] = 12'hB65;
w_real[104] = 12'h95A; w_imag[104] = 12'hB8F;
w_real[105] = 12'h93E; w_imag[105] = 12'hBB9;
w_real[106] = 12'h924; w_imag[106] = 12'hBE4;
w_real[107] = 12'h90B; w_imag[107] = 12'hC0F;
w_real[108] = 12'h8F2; w_imag[108] = 12'hC3B;
w_real[109] = 12'h8DB; w_imag[109] = 12'hC68;
w_real[110] = 12'h8C5; w_imag[110] = 12'hC95;
w_real[111] = 12'h8B0; w_imag[111] = 12'hCC3;
w_real[112] = 12'h89C; w_imag[112] = 12'hCF1;
w_real[113] = 12'h88A; w_imag[113] = 12'hD1F;
w_real[114] = 12'h878; w_imag[114] = 12'hD4F;
w_real[115] = 12'h868; w_imag[115] = 12'hD7E;
w_real[116] = 12'h859; w_imag[116] = 12'hDAE;
w_real[117] = 12'h84B; w_imag[117] = 12'hDDE;
w_real[118] = 12'h83E; w_imag[118] = 12'hE0F;
w_real[119] = 12'h832; w_imag[119] = 12'hE40;
w_real[120] = 12'h828; w_imag[120] = 12'hE71;
w_real[121] = 12'h81F; w_imag[121] = 12'hEA2;
w_real[122] = 12'h817; w_imag[122] = 12'hED4;
w_real[123] = 12'h810; w_imag[123] = 12'hF06;
w_real[124] = 12'h80A; w_imag[124] = 12'hF38;
w_real[125] = 12'h806; w_imag[125] = 12'hF6A;
w_real[126] = 12'h803; w_imag[126] = 12'hF9C;
w_real[127] = 12'h801; w_imag[127] = 12'hFCE;
w_real[128] = 12'h800; w_imag[128] = 12'h000;
w_real[129] = 12'h801; w_imag[129] = 12'h032;
w_real[130] = 12'h803; w_imag[130] = 12'h064;
w_real[131] = 12'h806; w_imag[131] = 12'h096;
w_real[132] = 12'h80A; w_imag[132] = 12'h0C8;
w_real[133] = 12'h810; w_imag[133] = 12'h0FA;
w_real[134] = 12'h817; w_imag[134] = 12'h12C;
w_real[135] = 12'h81F; w_imag[135] = 12'h15E;
w_real[136] = 12'h828; w_imag[136] = 12'h18F;
w_real[137] = 12'h832; w_imag[137] = 12'h1C0;
w_real[138] = 12'h83E; w_imag[138] = 12'h1F1;
w_real[139] = 12'h84B; w_imag[139] = 12'h222;
w_real[140] = 12'h859; w_imag[140] = 12'h252;
w_real[141] = 12'h868; w_imag[141] = 12'h282;
w_real[142] = 12'h878; w_imag[142] = 12'h2B1;
w_real[143] = 12'h88A; w_imag[143] = 12'h2E1;
w_real[144] = 12'h89C; w_imag[144] = 12'h30F;
w_real[145] = 12'h8B0; w_imag[145] = 12'h33D;
w_real[146] = 12'h8C5; w_imag[146] = 12'h36B;
w_real[147] = 12'h8DB; w_imag[147] = 12'h398;
w_real[148] = 12'h8F2; w_imag[148] = 12'h3C5;
w_real[149] = 12'h90B; w_imag[149] = 12'h3F1;
w_real[150] = 12'h924; w_imag[150] = 12'h41C;
w_real[151] = 12'h93E; w_imag[151] = 12'h447;
w_real[152] = 12'h95A; w_imag[152] = 12'h471;
w_real[153] = 12'h976; w_imag[153] = 12'h49B;
w_real[154] = 12'h994; w_imag[154] = 12'h4C3;
w_real[155] = 12'h9B2; w_imag[155] = 12'h4EB;
w_real[156] = 12'h9D1; w_imag[156] = 12'h513;
w_real[157] = 12'h9F2; w_imag[157] = 12'h539;
w_real[158] = 12'hA13; w_imag[158] = 12'h55F;
w_real[159] = 12'hA35; w_imag[159] = 12'h584;
w_real[160] = 12'hA58; w_imag[160] = 12'h5A8;
w_real[161] = 12'hA7C; w_imag[161] = 12'h5CB;
w_real[162] = 12'hAA1; w_imag[162] = 12'h5ED;
w_real[163] = 12'hAC7; w_imag[163] = 12'h60E;
w_real[164] = 12'hAED; w_imag[164] = 12'h62F;
w_real[165] = 12'hB15; w_imag[165] = 12'h64E;
w_real[166] = 12'hB3D; w_imag[166] = 12'h66C;
w_real[167] = 12'hB65; w_imag[167] = 12'h68A;
w_real[168] = 12'hB8F; w_imag[168] = 12'h6A6;
w_real[169] = 12'hBB9; w_imag[169] = 12'h6C2;
w_real[170] = 12'hBE4; w_imag[170] = 12'h6DC;
w_real[171] = 12'hC0F; w_imag[171] = 12'h6F5;
w_real[172] = 12'hC3B; w_imag[172] = 12'h70E;
w_real[173] = 12'hC68; w_imag[173] = 12'h725;
w_real[174] = 12'hC95; w_imag[174] = 12'h73B;
w_real[175] = 12'hCC3; w_imag[175] = 12'h750;
w_real[176] = 12'hCF1; w_imag[176] = 12'h764;
w_real[177] = 12'hD1F; w_imag[177] = 12'h776;
w_real[178] = 12'hD4F; w_imag[178] = 12'h788;
w_real[179] = 12'hD7E; w_imag[179] = 12'h798;
w_real[180] = 12'hDAE; w_imag[180] = 12'h7A7;
w_real[181] = 12'hDDE; w_imag[181] = 12'h7B5;
w_real[182] = 12'hE0F; w_imag[182] = 12'h7C2;
w_real[183] = 12'hE40; w_imag[183] = 12'h7CE;
w_real[184] = 12'hE71; w_imag[184] = 12'h7D8;
w_real[185] = 12'hEA2; w_imag[185] = 12'h7E1;
w_real[186] = 12'hED4; w_imag[186] = 12'h7E9;
w_real[187] = 12'hF06; w_imag[187] = 12'h7F0;
w_real[188] = 12'hF38; w_imag[188] = 12'h7F6;
w_real[189] = 12'hF6A; w_imag[189] = 12'h7FA;
w_real[190] = 12'hF9C; w_imag[190] = 12'h7FD;
w_real[191] = 12'hFCE; w_imag[191] = 12'h7FF;
w_real[192] = 12'h000; w_imag[192] = 12'h7FF;
w_real[193] = 12'h032; w_imag[193] = 12'h7FF;
w_real[194] = 12'h064; w_imag[194] = 12'h7FD;
w_real[195] = 12'h096; w_imag[195] = 12'h7FA;
w_real[196] = 12'h0C8; w_imag[196] = 12'h7F6;
w_real[197] = 12'h0FA; w_imag[197] = 12'h7F0;
w_real[198] = 12'h12C; w_imag[198] = 12'h7E9;
w_real[199] = 12'h15E; w_imag[199] = 12'h7E1;
w_real[200] = 12'h18F; w_imag[200] = 12'h7D8;
w_real[201] = 12'h1C0; w_imag[201] = 12'h7CE;
w_real[202] = 12'h1F1; w_imag[202] = 12'h7C2;
w_real[203] = 12'h222; w_imag[203] = 12'h7B5;
w_real[204] = 12'h252; w_imag[204] = 12'h7A7;
w_real[205] = 12'h282; w_imag[205] = 12'h798;
w_real[206] = 12'h2B1; w_imag[206] = 12'h788;
w_real[207] = 12'h2E1; w_imag[207] = 12'h776;
w_real[208] = 12'h30F; w_imag[208] = 12'h764;
w_real[209] = 12'h33D; w_imag[209] = 12'h750;
w_real[210] = 12'h36B; w_imag[210] = 12'h73B;
w_real[211] = 12'h398; w_imag[211] = 12'h725;
w_real[212] = 12'h3C5; w_imag[212] = 12'h70E;
w_real[213] = 12'h3F1; w_imag[213] = 12'h6F5;
w_real[214] = 12'h41C; w_imag[214] = 12'h6DC;
w_real[215] = 12'h447; w_imag[215] = 12'h6C2;
w_real[216] = 12'h471; w_imag[216] = 12'h6A6;
w_real[217] = 12'h49B; w_imag[217] = 12'h68A;
w_real[218] = 12'h4C3; w_imag[218] = 12'h66C;
w_real[219] = 12'h4EB; w_imag[219] = 12'h64E;
w_real[220] = 12'h513; w_imag[220] = 12'h62F;
w_real[221] = 12'h539; w_imag[221] = 12'h60E;
w_real[222] = 12'h55F; w_imag[222] = 12'h5ED;
w_real[223] = 12'h584; w_imag[223] = 12'h5CB;
w_real[224] = 12'h5A8; w_imag[224] = 12'h5A8;
w_real[225] = 12'h5CB; w_imag[225] = 12'h584;
w_real[226] = 12'h5ED; w_imag[226] = 12'h55F;
w_real[227] = 12'h60E; w_imag[227] = 12'h539;
w_real[228] = 12'h62F; w_imag[228] = 12'h513;
w_real[229] = 12'h64E; w_imag[229] = 12'h4EB;
w_real[230] = 12'h66C; w_imag[230] = 12'h4C3;
w_real[231] = 12'h68A; w_imag[231] = 12'h49B;
w_real[232] = 12'h6A6; w_imag[232] = 12'h471;
w_real[233] = 12'h6C2; w_imag[233] = 12'h447;
w_real[234] = 12'h6DC; w_imag[234] = 12'h41C;
w_real[235] = 12'h6F5; w_imag[235] = 12'h3F1;
w_real[236] = 12'h70E; w_imag[236] = 12'h3C5;
w_real[237] = 12'h725; w_imag[237] = 12'h398;
w_real[238] = 12'h73B; w_imag[238] = 12'h36B;
w_real[239] = 12'h750; w_imag[239] = 12'h33D;
w_real[240] = 12'h764; w_imag[240] = 12'h30F;
w_real[241] = 12'h776; w_imag[241] = 12'h2E1;
w_real[242] = 12'h788; w_imag[242] = 12'h2B1;
w_real[243] = 12'h798; w_imag[243] = 12'h282;
w_real[244] = 12'h7A7; w_imag[244] = 12'h252;
w_real[245] = 12'h7B5; w_imag[245] = 12'h222;
w_real[246] = 12'h7C2; w_imag[246] = 12'h1F1;
w_real[247] = 12'h7CE; w_imag[247] = 12'h1C0;
w_real[248] = 12'h7D8; w_imag[248] = 12'h18F;
w_real[249] = 12'h7E1; w_imag[249] = 12'h15E;
w_real[250] = 12'h7E9; w_imag[250] = 12'h12C;
w_real[251] = 12'h7F0; w_imag[251] = 12'h0FA;
w_real[252] = 12'h7F6; w_imag[252] = 12'h0C8;
w_real[253] = 12'h7FA; w_imag[253] = 12'h096;
w_real[254] = 12'h7FD; w_imag[254] = 12'h064;
w_real[255] = 12'h7FF; w_imag[255] = 12'h032;
