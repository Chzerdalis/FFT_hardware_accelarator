0 0
0 -14
2 -28
6 -43
14 -74
20 -83
43 -142
43 -120
62 -151
96 -203
152 -286
459 -766
706 -1057
107 -145
986 -1202
525 -579
667 -667
800 -725
-314 257
-653 484
-425 284
-321 192
-151 80
-179 84
-320 132
-411 147
-332 100
-293 73
-299 59
-290 43
-283 27
-278 13
-282 0
-278 -13
-283 -27
-290 -43
-299 -59
-293 -73
-332 -100
-411 -147
-320 -132
-179 -84
-151 -80
-321 -192
-425 -284
-653 -484
-314 -257
800 725
667 667
525 579
986 1202
107 145
706 1057
459 766
152 286
96 203
62 151
43 120
43 142
20 83
14 74
6 43
2 28
0 14
